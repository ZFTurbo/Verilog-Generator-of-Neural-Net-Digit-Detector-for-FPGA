module database(clk,datata,re,address,we,dp,address_p);

parameter SIZE=0;

input clk;
output reg signed [SIZE-1:0] datata;
input re,we;
input [12:0] address;
input signed [SIZE-1:0] dp;
input [12:0] address_p;

reg signed [SIZE-1:0] storage [5459:0];

initial begin

storage[0] =  12'b0;
storage[1] =  12'b0;
storage[2] =  12'b0;
storage[3] =  12'b0;
storage[4] =  12'b0;
storage[5] =  12'b0;
storage[6] =  12'b0;
storage[7] =  12'b0;
storage[8] =  12'b0;
storage[9] =  12'b0;
storage[10] =  12'b0;
storage[11] =  12'b0;
storage[12] =  12'b0;
storage[13] =  12'b0;
storage[14] =  12'b0;
storage[15] =  12'b0;
storage[16] =  12'b0;
storage[17] =  12'b0;
storage[18] =  12'b0;
storage[19] =  12'b0;
storage[20] =  12'b0;
storage[21] =  12'b0;
storage[22] =  12'b0;
storage[23] =  12'b0;
storage[24] =  12'b0;
storage[25] =  12'b0;
storage[26] =  12'b0;
storage[27] =  12'b0;
storage[28] =  12'b0;
storage[29] =  12'b0;
storage[30] =  12'b0;
storage[31] =  12'b0;
storage[32] =  12'b0;
storage[33] =  12'b0;
storage[34] =  12'b0;
storage[35] =  12'b0;
storage[36] =  12'b0;
storage[37] =  12'b0;
storage[38] =  12'b0;
storage[39] =  12'b0;
storage[40] =  12'b0;
storage[41] =  12'b0;
storage[42] =  12'b0;
storage[43] =  12'b0;
storage[44] =  12'b0;
storage[45] =  12'b0;
storage[46] =  12'b0;
storage[47] =  12'b0;
storage[48] =  12'b0;
storage[49] =  12'b0;
storage[50] =  12'b0;
storage[51] =  12'b0;
storage[52] =  12'b0;
storage[53] =  12'b0;
storage[54] =  12'b0;
storage[55] =  12'b0;
storage[56] =  12'b0;
storage[57] =  12'b0;
storage[58] =  12'b0;
storage[59] =  12'b0;
storage[60] =  12'b0;
storage[61] =  12'b0;
storage[62] =  12'b0;
storage[63] =  12'b0;
storage[64] =  12'b0;
storage[65] =  12'b0;
storage[66] =  12'b0;
storage[67] =  12'b0;
storage[68] =  12'b0;
storage[69] =  12'b0;
storage[70] =  12'b0;
storage[71] =  12'b0;
storage[72] =  12'b0;
storage[73] =  12'b0;
storage[74] =  12'b0;
storage[75] =  12'b0;
storage[76] =  12'b0;
storage[77] =  12'b0;
storage[78] =  12'b0;
storage[79] =  12'b0;
storage[80] =  12'b0;
storage[81] =  12'b0;
storage[82] =  12'b0;
storage[83] =  12'b0;
storage[84] =  12'b0;
storage[85] =  12'b0;
storage[86] =  12'b0;
storage[87] =  12'b0;
storage[88] =  12'b0;
storage[89] =  12'b0;
storage[90] =  12'b0;
storage[91] =  12'b0;
storage[92] =  12'b0;
storage[93] =  12'b0;
storage[94] =  12'b0;
storage[95] =  12'b0;
storage[96] =  12'b0;
storage[97] =  12'b0;
storage[98] =  12'b0;
storage[99] =  12'b0;
storage[100] =  12'b0;
storage[101] =  12'b0;
storage[102] =  12'b0;
storage[103] =  12'b0;
storage[104] =  12'b0;
storage[105] =  12'b0;
storage[106] =  12'b0;
storage[107] =  12'b0;
storage[108] =  12'b0;
storage[109] =  12'b0;
storage[110] =  12'b0;
storage[111] =  12'b0;
storage[112] =  12'b0;
storage[113] =  12'b0;
storage[114] =  12'b0;
storage[115] =  12'b0;
storage[116] =  12'b0;
storage[117] =  12'b0;
storage[118] =  12'b0;
storage[119] =  12'b0;
storage[120] =  12'b0;
storage[121] =  12'b0;
storage[122] =  12'b0;
storage[123] =  12'b0;
storage[124] =  12'b0;
storage[125] =  12'b0;
storage[126] =  12'b0;
storage[127] =  12'b0;
storage[128] =  12'b0;
storage[129] =  12'b0;
storage[130] =  12'b0;
storage[131] =  12'b0;
storage[132] =  12'b0;
storage[133] =  12'b0;
storage[134] =  12'b0;
storage[135] =  12'b0;
storage[136] =  12'b0;
storage[137] =  12'b0;
storage[138] =  12'b0;
storage[139] =  12'b0;
storage[140] =  12'b0;
storage[141] =  12'b0;
storage[142] =  12'b0;
storage[143] =  12'b0;
storage[144] =  12'b0;
storage[145] =  12'b0;
storage[146] =  12'b0;
storage[147] =  12'b0;
storage[148] =  12'b0;
storage[149] =  12'b0;
storage[150] =  12'b0;
storage[151] =  12'b0;
storage[152] =  12'b0;
storage[153] =  12'b0;
storage[154] =  12'b0;
storage[155] =  12'b0;
storage[156] =  12'b0;
storage[157] =  12'b0;
storage[158] =  12'b0;
storage[159] =  12'b0;
storage[160] =  12'b0;
storage[161] =  12'b0;
storage[162] =  12'b0;
storage[163] =  12'b0;
storage[164] =  12'b0;
storage[165] =  12'b0;
storage[166] =  12'b0;
storage[167] =  12'b0;
storage[168] =  12'b0;
storage[169] =  12'b0;
storage[170] =  12'b0;
storage[171] =  12'b0;
storage[172] =  12'b0;
storage[173] =  12'b0;
storage[174] =  12'b0;
storage[175] =  12'b0;
storage[176] =  12'b0;
storage[177] =  12'b0;
storage[178] =  12'b0;
storage[179] =  12'b0;
storage[180] =  12'b0;
storage[181] =  12'b0;
storage[182] =  12'b0;
storage[183] =  12'b0;
storage[184] =  12'b0;
storage[185] =  12'b0;
storage[186] =  12'b0;
storage[187] =  12'b0;
storage[188] =  12'b0;
storage[189] =  12'b0;
storage[190] =  12'b0;
storage[191] =  12'b0;
storage[192] =  12'b0;
storage[193] =  12'b0;
storage[194] =  12'b0;
storage[195] =  12'b0;
storage[196] =  12'b0;
storage[197] =  12'b0;
storage[198] =  12'b0;
storage[199] =  12'b0;
storage[200] =  12'b0;
storage[201] =  12'b0;
storage[202] =  12'b0;
storage[203] =  12'b0;
storage[204] =  12'b0;
storage[205] =  12'b0;
storage[206] =  12'b0;
storage[207] =  12'b0;
storage[208] =  12'b0;
storage[209] =  12'b0;
storage[210] =  12'b0;
storage[211] =  12'b0;
storage[212] =  12'b0;
storage[213] =  12'b0;
storage[214] =  12'b0;
storage[215] =  12'b0;
storage[216] =  12'b0;
storage[217] =  12'b0;
storage[218] =  12'b0;
storage[219] =  12'b0;
storage[220] =  12'b0;
storage[221] =  12'b0;
storage[222] =  12'b0;
storage[223] =  12'b0;
storage[224] =  12'b0;
storage[225] =  12'b0;
storage[226] =  12'b0;
storage[227] =  12'b0;
storage[228] =  12'b0;
storage[229] =  12'b0;
storage[230] =  12'b0;
storage[231] =  12'b0;
storage[232] =  12'b0;
storage[233] =  12'b0;
storage[234] =  12'b0;
storage[235] =  12'b0;
storage[236] =  12'b0;
storage[237] =  12'b0;
storage[238] =  12'b0;
storage[239] =  12'b0;
storage[240] =  12'b0;
storage[241] =  12'b0;
storage[242] =  12'b0;
storage[243] =  12'b0;
storage[244] =  12'b0;
storage[245] =  12'b0;
storage[246] =  12'b0;
storage[247] =  12'b0;
storage[248] =  12'b0;
storage[249] =  12'b0;
storage[250] =  12'b0;
storage[251] =  12'b0;
storage[252] =  12'b0;
storage[253] =  12'b0;
storage[254] =  12'b0;
storage[255] =  12'b0;
storage[256] =  12'b0;
storage[257] =  12'b0;
storage[258] =  12'b0;
storage[259] =  12'b0;
storage[260] =  12'b0;
storage[261] =  12'b0;
storage[262] =  12'b0;
storage[263] =  12'b0;
storage[264] =  12'b0;
storage[265] =  12'b0;
storage[266] =  12'b0;
storage[267] =  12'b0;
storage[268] =  12'b0;
storage[269] =  12'b0;
storage[270] =  12'b0;
storage[271] =  12'b0;
storage[272] =  12'b0;
storage[273] =  12'b0;
storage[274] =  12'b0;
storage[275] =  12'b0;
storage[276] =  12'b0;
storage[277] =  12'b0;
storage[278] =  12'b0;
storage[279] =  12'b0;
storage[280] =  12'b0;
storage[281] =  12'b0;
storage[282] =  12'b0;
storage[283] =  12'b0;
storage[284] =  12'b0;
storage[285] =  12'b0;
storage[286] =  12'b0;
storage[287] =  12'b0;
storage[288] =  12'b0;
storage[289] =  12'b0;
storage[290] =  12'b0;
storage[291] =  12'b0;
storage[292] =  12'b0;
storage[293] =  12'b0;
storage[294] =  12'b0;
storage[295] =  12'b0;
storage[296] =  12'b0;
storage[297] =  12'b0;
storage[298] =  12'b0;
storage[299] =  12'b0;
storage[300] =  12'b0;
storage[301] =  12'b0;
storage[302] =  12'b0;
storage[303] =  12'b0;
storage[304] =  12'b0;
storage[305] =  12'b0;
storage[306] =  12'b0;
storage[307] =  12'b0;
storage[308] =  12'b0;
storage[309] =  12'b0;
storage[310] =  12'b0;
storage[311] =  12'b0;
storage[312] =  12'b0;
storage[313] =  12'b0;
storage[314] =  12'b0;
storage[315] =  12'b0;
storage[316] =  12'b0;
storage[317] =  12'b0;
storage[318] =  12'b0;
storage[319] =  12'b0;
storage[320] =  12'b0;
storage[321] =  12'b0;
storage[322] =  12'b0;
storage[323] =  12'b0;
storage[324] =  12'b0;
storage[325] =  12'b0;
storage[326] =  12'b0;
storage[327] =  12'b0;
storage[328] =  12'b0;
storage[329] =  12'b0;
storage[330] =  12'b0;
storage[331] =  12'b0;
storage[332] =  12'b0;
storage[333] =  12'b0;
storage[334] =  12'b0;
storage[335] =  12'b0;
storage[336] =  12'b0;
storage[337] =  12'b0;
storage[338] =  12'b0;
storage[339] =  12'b0;
storage[340] =  12'b0;
storage[341] =  12'b0;
storage[342] =  12'b0;
storage[343] =  12'b0;
storage[344] =  12'b0;
storage[345] =  12'b0;
storage[346] =  12'b0;
storage[347] =  12'b0;
storage[348] =  12'b0;
storage[349] =  12'b0;
storage[350] =  12'b0;
storage[351] =  12'b0;
storage[352] =  12'b0;
storage[353] =  12'b0;
storage[354] =  12'b0;
storage[355] =  12'b0;
storage[356] =  12'b0;
storage[357] =  12'b0;
storage[358] =  12'b0;
storage[359] =  12'b0;
storage[360] =  12'b0;
storage[361] =  12'b0;
storage[362] =  12'b0;
storage[363] =  12'b0;
storage[364] =  12'b0;
storage[365] =  12'b0;
storage[366] =  12'b0;
storage[367] =  12'b0;
storage[368] =  12'b0;
storage[369] =  12'b0;
storage[370] =  12'b0;
storage[371] =  12'b0;
storage[372] =  12'b0;
storage[373] =  12'b0;
storage[374] =  12'b0;
storage[375] =  12'b0;
storage[376] =  12'b0;
storage[377] =  12'b0;
storage[378] =  12'b0;
storage[379] =  12'b0;
storage[380] =  12'b0;
storage[381] =  12'b0;
storage[382] =  12'b0;
storage[383] =  12'b0;
storage[384] =  12'b0;
storage[385] =  12'b0;
storage[386] =  12'b0;
storage[387] =  12'b0;
storage[388] =  12'b0;
storage[389] =  12'b0;
storage[390] =  12'b0;
storage[391] =  12'b0;
storage[392] =  12'b0;
storage[393] =  12'b0;
storage[394] =  12'b0;
storage[395] =  12'b0;
storage[396] =  12'b0;
storage[397] =  12'b0;
storage[398] =  12'b0;
storage[399] =  12'b0;
storage[400] =  12'b0;
storage[401] =  12'b0;
storage[402] =  12'b0;
storage[403] =  12'b0;
storage[404] =  12'b0;
storage[405] =  12'b0;
storage[406] =  12'b0;
storage[407] =  12'b0;
storage[408] =  12'b0;
storage[409] =  12'b0;
storage[410] =  12'b0;
storage[411] =  12'b0;
storage[412] =  12'b0;
storage[413] =  12'b0;
storage[414] =  12'b0;
storage[415] =  12'b0;
storage[416] =  12'b0;
storage[417] =  12'b0;
storage[418] =  12'b0;
storage[419] =  12'b0;
storage[420] =  12'b0;
storage[421] =  12'b0;
storage[422] =  12'b0;
storage[423] =  12'b0;
storage[424] =  12'b0;
storage[425] =  12'b0;
storage[426] =  12'b0;
storage[427] =  12'b0;
storage[428] =  12'b0;
storage[429] =  12'b0;
storage[430] =  12'b0;
storage[431] =  12'b0;
storage[432] =  12'b0;
storage[433] =  12'b0;
storage[434] =  12'b0;
storage[435] =  12'b0;
storage[436] =  12'b0;
storage[437] =  12'b0;
storage[438] =  12'b0;
storage[439] =  12'b0;
storage[440] =  12'b0;
storage[441] =  12'b0;
storage[442] =  12'b0;
storage[443] =  12'b0;
storage[444] =  12'b0;
storage[445] =  12'b0;
storage[446] =  12'b0;
storage[447] =  12'b0;
storage[448] =  12'b0;
storage[449] =  12'b0;
storage[450] =  12'b0;
storage[451] =  12'b0;
storage[452] =  12'b0;
storage[453] =  12'b0;
storage[454] =  12'b0;
storage[455] =  12'b0;
storage[456] =  12'b0;
storage[457] =  12'b0;
storage[458] =  12'b0;
storage[459] =  12'b0;
storage[460] =  12'b0;
storage[461] =  12'b0;
storage[462] =  12'b0;
storage[463] =  12'b0;
storage[464] =  12'b0;
storage[465] =  12'b0;
storage[466] =  12'b0;
storage[467] =  12'b0;
storage[468] =  12'b0;
storage[469] =  12'b0;
storage[470] =  12'b0;
storage[471] =  12'b0;
storage[472] =  12'b0;
storage[473] =  12'b0;
storage[474] =  12'b0;
storage[475] =  12'b0;
storage[476] =  12'b0;
storage[477] =  12'b0;
storage[478] =  12'b0;
storage[479] =  12'b0;
storage[480] =  12'b0;
storage[481] =  12'b0;
storage[482] =  12'b0;
storage[483] =  12'b0;
storage[484] =  12'b0;
storage[485] =  12'b0;
storage[486] =  12'b0;
storage[487] =  12'b0;
storage[488] =  12'b0;
storage[489] =  12'b0;
storage[490] =  12'b0;
storage[491] =  12'b0;
storage[492] =  12'b0;
storage[493] =  12'b0;
storage[494] =  12'b0;
storage[495] =  12'b0;
storage[496] =  12'b0;
storage[497] =  12'b0;
storage[498] =  12'b0;
storage[499] =  12'b0;
storage[500] =  12'b0;
storage[501] =  12'b0;
storage[502] =  12'b0;
storage[503] =  12'b0;
storage[504] =  12'b0;
storage[505] =  12'b0;
storage[506] =  12'b0;
storage[507] =  12'b0;
storage[508] =  12'b0;
storage[509] =  12'b0;
storage[510] =  12'b0;
storage[511] =  12'b0;
storage[512] =  12'b0;
storage[513] =  12'b0;
storage[514] =  12'b0;
storage[515] =  12'b0;
storage[516] =  12'b0;
storage[517] =  12'b0;
storage[518] =  12'b0;
storage[519] =  12'b0;
storage[520] =  12'b0;
storage[521] =  12'b0;
storage[522] =  12'b0;
storage[523] =  12'b0;
storage[524] =  12'b0;
storage[525] =  12'b0;
storage[526] =  12'b0;
storage[527] =  12'b0;
storage[528] =  12'b0;
storage[529] =  12'b0;
storage[530] =  12'b0;
storage[531] =  12'b0;
storage[532] =  12'b0;
storage[533] =  12'b0;
storage[534] =  12'b0;
storage[535] =  12'b0;
storage[536] =  12'b0;
storage[537] =  12'b0;
storage[538] =  12'b0;
storage[539] =  12'b0;
storage[540] =  12'b0;
storage[541] =  12'b0;
storage[542] =  12'b0;
storage[543] =  12'b0;
storage[544] =  12'b0;
storage[545] =  12'b0;
storage[546] =  12'b0;
storage[547] =  12'b0;
storage[548] =  12'b0;
storage[549] =  12'b0;
storage[550] =  12'b0;
storage[551] =  12'b0;
storage[552] =  12'b0;
storage[553] =  12'b0;
storage[554] =  12'b0;
storage[555] =  12'b0;
storage[556] =  12'b0;
storage[557] =  12'b0;
storage[558] =  12'b0;
storage[559] =  12'b0;
storage[560] =  12'b0;
storage[561] =  12'b0;
storage[562] =  12'b0;
storage[563] =  12'b0;
storage[564] =  12'b0;
storage[565] =  12'b0;
storage[566] =  12'b0;
storage[567] =  12'b0;
storage[568] =  12'b0;
storage[569] =  12'b0;
storage[570] =  12'b0;
storage[571] =  12'b0;
storage[572] =  12'b0;
storage[573] =  12'b0;
storage[574] =  12'b0;
storage[575] =  12'b0;
storage[576] =  12'b0;
storage[577] =  12'b0;
storage[578] =  12'b0;
storage[579] =  12'b0;
storage[580] =  12'b0;
storage[581] =  12'b0;
storage[582] =  12'b0;
storage[583] =  12'b0;
storage[584] =  12'b0;
storage[585] =  12'b0;
storage[586] =  12'b0;
storage[587] =  12'b0;
storage[588] =  12'b0;
storage[589] =  12'b0;
storage[590] =  12'b0;
storage[591] =  12'b0;
storage[592] =  12'b0;
storage[593] =  12'b0;
storage[594] =  12'b0;
storage[595] =  12'b0;
storage[596] =  12'b0;
storage[597] =  12'b0;
storage[598] =  12'b0;
storage[599] =  12'b0;
storage[600] =  12'b0;
storage[601] =  12'b0;
storage[602] =  12'b0;
storage[603] =  12'b0;
storage[604] =  12'b0;
storage[605] =  12'b0;
storage[606] =  12'b0;
storage[607] =  12'b0;
storage[608] =  12'b0;
storage[609] =  12'b0;
storage[610] =  12'b0;
storage[611] =  12'b0;
storage[612] =  12'b0;
storage[613] =  12'b0;
storage[614] =  12'b0;
storage[615] =  12'b0;
storage[616] =  12'b0;
storage[617] =  12'b0;
storage[618] =  12'b0;
storage[619] =  12'b0;
storage[620] =  12'b0;
storage[621] =  12'b0;
storage[622] =  12'b0;
storage[623] =  12'b0;
storage[624] =  12'b0;
storage[625] =  12'b0;
storage[626] =  12'b0;
storage[627] =  12'b0;
storage[628] =  12'b0;
storage[629] =  12'b0;
storage[630] =  12'b0;
storage[631] =  12'b0;
storage[632] =  12'b0;
storage[633] =  12'b0;
storage[634] =  12'b0;
storage[635] =  12'b0;
storage[636] =  12'b0;
storage[637] =  12'b0;
storage[638] =  12'b0;
storage[639] =  12'b0;
storage[640] =  12'b0;
storage[641] =  12'b0;
storage[642] =  12'b0;
storage[643] =  12'b0;
storage[644] =  12'b0;
storage[645] =  12'b0;
storage[646] =  12'b0;
storage[647] =  12'b0;
storage[648] =  12'b0;
storage[649] =  12'b0;
storage[650] =  12'b0;
storage[651] =  12'b0;
storage[652] =  12'b0;
storage[653] =  12'b0;
storage[654] =  12'b0;
storage[655] =  12'b0;
storage[656] =  12'b0;
storage[657] =  12'b0;
storage[658] =  12'b0;
storage[659] =  12'b0;
storage[660] =  12'b0;
storage[661] =  12'b0;
storage[662] =  12'b0;
storage[663] =  12'b0;
storage[664] =  12'b0;
storage[665] =  12'b0;
storage[666] =  12'b0;
storage[667] =  12'b0;
storage[668] =  12'b0;
storage[669] =  12'b0;
storage[670] =  12'b0;
storage[671] =  12'b0;
storage[672] =  12'b0;
storage[673] =  12'b0;
storage[674] =  12'b0;
storage[675] =  12'b0;
storage[676] =  12'b0;
storage[677] =  12'b0;
storage[678] =  12'b0;
storage[679] =  12'b0;
storage[680] =  12'b0;
storage[681] =  12'b0;
storage[682] =  12'b0;
storage[683] =  12'b0;
storage[684] =  12'b0;
storage[685] =  12'b0;
storage[686] =  12'b0;
storage[687] =  12'b0;
storage[688] =  12'b0;
storage[689] =  12'b0;
storage[690] =  12'b0;
storage[691] =  12'b0;
storage[692] =  12'b0;
storage[693] =  12'b0;
storage[694] =  12'b0;
storage[695] =  12'b0;
storage[696] =  12'b0;
storage[697] =  12'b0;
storage[698] =  12'b0;
storage[699] =  12'b0;
storage[700] =  12'b0;
storage[701] =  12'b0;
storage[702] =  12'b0;
storage[703] =  12'b0;
storage[704] =  12'b0;
storage[705] =  12'b0;
storage[706] =  12'b0;
storage[707] =  12'b0;
storage[708] =  12'b0;
storage[709] =  12'b0;
storage[710] =  12'b0;
storage[711] =  12'b0;
storage[712] =  12'b0;
storage[713] =  12'b0;
storage[714] =  12'b0;
storage[715] =  12'b0;
storage[716] =  12'b0;
storage[717] =  12'b0;
storage[718] =  12'b0;
storage[719] =  12'b0;
storage[720] =  12'b0;
storage[721] =  12'b0;
storage[722] =  12'b0;
storage[723] =  12'b0;
storage[724] =  12'b0;
storage[725] =  12'b0;
storage[726] =  12'b0;
storage[727] =  12'b0;
storage[728] =  12'b0;
storage[729] =  12'b0;
storage[730] =  12'b0;
storage[731] =  12'b0;
storage[732] =  12'b0;
storage[733] =  12'b0;
storage[734] =  12'b0;
storage[735] =  12'b0;
storage[736] =  12'b0;
storage[737] =  12'b0;
storage[738] =  12'b0;
storage[739] =  12'b0;
storage[740] =  12'b0;
storage[741] =  12'b0;
storage[742] =  12'b0;
storage[743] =  12'b0;
storage[744] =  12'b0;
storage[745] =  12'b0;
storage[746] =  12'b0;
storage[747] =  12'b0;
storage[748] =  12'b0;
storage[749] =  12'b0;
storage[750] =  12'b0;
storage[751] =  12'b0;
storage[752] =  12'b0;
storage[753] =  12'b0;
storage[754] =  12'b0;
storage[755] =  12'b0;
storage[756] =  12'b0;
storage[757] =  12'b0;
storage[758] =  12'b0;
storage[759] =  12'b0;
storage[760] =  12'b0;
storage[761] =  12'b0;
storage[762] =  12'b0;
storage[763] =  12'b0;
storage[764] =  12'b0;
storage[765] =  12'b0;
storage[766] =  12'b0;
storage[767] =  12'b0;
storage[768] =  12'b0;
storage[769] =  12'b0;
storage[770] =  12'b0;
storage[771] =  12'b0;
storage[772] =  12'b0;
storage[773] =  12'b0;
storage[774] =  12'b0;
storage[775] =  12'b0;
storage[776] =  12'b0;
storage[777] =  12'b0;
storage[778] =  12'b0;
storage[779] =  12'b0;
storage[780] =  12'b0;
storage[781] =  12'b0;
storage[782] =  12'b0;
storage[783] =  12'b0;
storage[784] =  12'b000100101000; // 296
storage[785] =  12'b001001111010; // 634
storage[786] = -12'b000011010111; // -215
storage[787] = -12'b000001010010; // -82
storage[788] = -12'b000000110101; // -53
storage[789] = -12'b000000110111; // -55
storage[790] = -12'b000110000011; // -387
storage[791] =  12'b000101010111; // 343
storage[792] = -12'b000110000001; // -385
storage[793] = -12'b000010101110; // -174
storage[794] = -12'b000001110111; // -119
storage[795] =  12'b001000100000; // 544
storage[796] = -12'b000010110110; // -182
storage[797] = -12'b000001001001; // -73
storage[798] =  12'b000111000111; // 455
storage[799] = -12'b000011101001; // -233
storage[800] = -12'b000101010000; // -336
storage[801] =  12'b000011111010; // 250
storage[802] =  12'b000001100100; // 100
storage[803] = -12'b000100110101; // -309
storage[804] =  12'b000000010011; // 19
storage[805] = -12'b000100000000; // -256
storage[806] = -12'b000011000001; // -193
storage[807] = -12'b000010110011; // -179
storage[808] =  12'b000110011101; // 413
storage[809] =  12'b000110011001; // 409
storage[810] =  12'b000010011000; // 152
storage[811] =  12'b000010001110; // 142
storage[812] =  12'b000100000110; // 262
storage[813] =  12'b000100101001; // 297
storage[814] =  12'b000001011011; // 91
storage[815] =  12'b000111011100; // 476
storage[816] =  12'b000000101100; // 44
storage[817] =  12'b000100000101; // 261
storage[818] =  12'b000100101000; // 296
storage[819] = -12'b000010001100; // -140
storage[820] =  12'b000010001100; // 140
storage[821] =  12'b000011010100; // 212
storage[822] =  12'b000001111110; // 126
storage[823] = -12'b000010011111; // -159
storage[824] = -12'b001011111011; // -763
storage[825] = -12'b000111111001; // -505
storage[826] = -12'b000111011010; // -474
storage[827] = -12'b001100010100; // -788
storage[828] = -12'b000100001000; // -264
storage[829] = -12'b000100110100; // -308
storage[830] = -12'b000001000110; // -70
storage[831] = -12'b000001100101; // -101
storage[832] =  12'b000000000111; // 7
storage[833] = -12'b000001111000; // -120
storage[834] = -12'b000101001000; // -328
storage[835] =  12'b000011011010; // 218
storage[836] =  12'b000010011000; // 152
storage[837] = -12'b000000000011; // -3
storage[838] =  12'b000000100011; // 35
storage[839] =  12'b000100101010; // 298
storage[840] =  12'b000010100011; // 163
storage[841] =  12'b000001100010; // 98
storage[842] =  12'b000001001111; // 79
storage[843] =  12'b000111010011; // 467
storage[844] =  12'b000011100011; // 227
storage[845] =  12'b000011100111; // 231
storage[846] =  12'b000011001110; // 206
storage[847] =  12'b000010001000; // 136
storage[848] = -12'b000001000011; // -67
storage[849] =  12'b000000101010; // 42
storage[850] = -12'b000010011001; // -153
storage[851] =  12'b000000000100; // 4
storage[852] = -12'b000001100011; // -99
storage[853] = -12'b000011110101; // -245
storage[854] =  12'b000001001011; // 75
storage[855] =  12'b000011000011; // 195
storage[856] =  12'b000001110010; // 114
storage[857] = -12'b000110111001; // -441
storage[858] =  12'b000000101101; // 45
storage[859] = -12'b000010001101; // -141
storage[860] = -12'b000110000101; // -389
storage[861] =  12'b000100001101; // 269
storage[862] =  12'b000110001010; // 394
storage[863] = -12'b000001011000; // -88
storage[864] =  12'b000000010111; // 23
storage[865] = -12'b000101010110; // -342
storage[866] = -12'b000110011011; // -411
storage[867] =  12'b000001010100; // 84
storage[868] = -12'b000110010101; // -405
storage[869] = -12'b001001111110; // -638
storage[870] =  12'b000000111110; // 62
storage[871] = -12'b001010100101; // -677
storage[872] = -12'b001001101011; // -619
storage[873] = -12'b000011011111; // -223
storage[874] =  12'b000111001010; // 458
storage[875] =  12'b000101000000; // 320
storage[876] =  12'b000000100100; // 36
storage[877] =  12'b000100001001; // 265
storage[878] = -12'b000010010100; // -148
storage[879] =  12'b000000111010; // 58
storage[880] =  12'b000100101100; // 300
storage[881] = -12'b000001001001; // -73
storage[882] = -12'b000001011111; // -95
storage[883] =  12'b000100011100; // 284
storage[884] = -12'b000001101011; // -107
storage[885] = -12'b000010011110; // -158
storage[886] =  12'b000000001000; // 8
storage[887] = -12'b000000010011; // -19
storage[888] =  12'b000000011110; // 30
storage[889] =  12'b000100101101; // 301
storage[890] = -12'b000010010000; // -144
storage[891] = -12'b000011011100; // -220
storage[892] =  12'b000100001101; // 269
storage[893] = -12'b000011001001; // -201
storage[894] =  12'b000011100010; // 226
storage[895] =  12'b000000110000; // 48
storage[896] =  12'b000000001010; // 10
storage[897] =  12'b000110101101; // 429
storage[898] =  12'b000010100101; // 165
storage[899] =  12'b000010001110; // 142
storage[900] =  12'b000110100111; // 423
storage[901] = -12'b000010111001; // -185
storage[902] = -12'b000100001111; // -271
storage[903] = -12'b000011000111; // -199
storage[904] = -12'b000001001101; // -77
storage[905] = -12'b001001010100; // -596
storage[906] = -12'b000000010111; // -23
storage[907] =  12'b000111100000; // 480
storage[908] = -12'b000001010110; // -86
storage[909] =  12'b000001111000; // 120
storage[910] = -12'b000011000011; // -195
storage[911] = -12'b000001111111; // -127
storage[912] = -12'b000110110000; // -432
storage[913] =  12'b000001011101; // 93
storage[914] = -12'b000101001100; // -332
storage[915] = -12'b000100100111; // -295
storage[916] = -12'b000111010011; // -467
storage[917] = -12'b000100111010; // -314
storage[918] = -12'b000100111001; // -313
storage[919] = -12'b000001011100; // -92
storage[920] = -12'b000000100000; // -32
storage[921] = -12'b000000000101; // -5
storage[922] =  12'b000011010111; // 215
storage[923] =  12'b000001110101; // 117
storage[924] =  12'b000010110010; // 178
storage[925] =  12'b000000100001; // 33
storage[926] =  12'b000010001001; // 137
storage[927] =  12'b000000000111; // 7
storage[928] = -12'b000001100100; // -100
storage[929] = -12'b001010000011; // -643
storage[930] =  12'b000101010000; // 336
storage[931] = -12'b000011001010; // -202
storage[932] = -12'b000111101001; // -489
storage[933] = -12'b000010110100; // -180
storage[934] = -12'b000110001010; // -394
storage[935] = -12'b001000010100; // -532
storage[936] =  12'b000011111110; // 254
storage[937] =  12'b000010100101; // 165
storage[938] =  12'b000010100110; // 166
storage[939] =  12'b000010001111; // 143
storage[940] =  12'b000011110111; // 247
storage[941] =  12'b000100101011; // 299
storage[942] =  12'b000100000111; // 263
storage[943] =  12'b000100000101; // 261
storage[944] =  12'b000010001111; // 143
storage[945] =  12'b000011100110; // 230
storage[946] = -12'b000101010001; // -337
storage[947] = -12'b000000111000; // -56
storage[948] =  12'b000100001000; // 264
storage[949] = -12'b000010110100; // -180
storage[950] = -12'b001001000011; // -579
storage[951] = -12'b000011000100; // -196
storage[952] = -12'b000000110011; // -51
storage[953] = -12'b000011111111; // -255
storage[954] = -12'b000010110100; // -180
storage[955] =  12'b000010011111; // 159
storage[956] = -12'b000010010111; // -151
storage[957] = -12'b000000010011; // -19
storage[958] = -12'b000010110010; // -178
storage[959] = -12'b000000110111; // -55
storage[960] =  12'b000001001001; // 73
storage[961] =  12'b000001110110; // 118
storage[962] = -12'b000000110111; // -55
storage[963] =  12'b000010010111; // 151
storage[964] =  12'b000000101010; // 42
storage[965] = -12'b000110110111; // -439
storage[966] = -12'b011101000110; // -1862
storage[967] = -12'b000111111011; // -507
storage[968] = -12'b010100100000; // -1312
storage[969] = -12'b010010111001; // -1209
storage[970] = -12'b001000001111; // -527
storage[971] = -12'b001010101011; // -683
storage[972] = -12'b001001100001; // -609
storage[973] = -12'b000000100010; // -34
storage[974] = -12'b000011100011; // -227
storage[975] = -12'b000001000110; // -70
storage[976] =  12'b000001111001; // 121
storage[977] = -12'b000011111000; // -248
storage[978] =  12'b000011000110; // 198
storage[979] = -12'b000110001001; // -393
storage[980] =  12'b000100011111; // 287
storage[981] =  12'b001001110111; // 631
storage[982] = -12'b000011001011; // -203
storage[983] =  12'b000100111110; // 318
storage[984] = -12'b000101000111; // -327
storage[985] =  12'b000011000000; // 192
storage[986] =  12'b001000000111; // 519
storage[987] = -12'b000001011100; // -92
storage[988] =  12'b000100010000; // 272
storage[989] =  12'b000111101011; // 491
storage[990] = -12'b000011001000; // -200
storage[991] = -12'b000010111101; // -189
storage[992] =  12'b000001111010; // 122
storage[993] = -12'b000111111010; // -506
storage[994] = -12'b001000101100; // -556
storage[995] = -12'b001000100100; // -548
storage[996] = -12'b000110011001; // -409
storage[997] = -12'b000110101010; // -426
storage[998] = -12'b000100000110; // -262
storage[999] = -12'b000000100101; // -37
storage[1000] =  12'b000101101111; // 367
storage[1001] = -12'b000101100010; // -354
storage[1002] = -12'b001101101001; // -873
storage[1003] = -12'b001010110000; // -688
storage[1004] = -12'b010000001100; // -1036
storage[1005] = -12'b001010100011; // -675
storage[1006] = -12'b000000111111; // -63
storage[1007] =  12'b000001000001; // 65
storage[1008] =  12'b000011000111; // 199
storage[1009] = -12'b000101101001; // -361
storage[1010] =  12'b000011001100; // 204
storage[1011] =  12'b001001001010; // 586
storage[1012] = -12'b000110010011; // -403
storage[1013] = -12'b000001111001; // -121
storage[1014] =  12'b001000010100; // 532
storage[1015] = -12'b000000011000; // -24
storage[1016] =  12'b000010100001; // 161
storage[1017] =  12'b000000000001; // 1
storage[1018] = -12'b000000011111; // -31
storage[1019] = -12'b000101000000; // -320
storage[1020] = -12'b000010101000; // -168
storage[1021] =  12'b000110011101; // 413
storage[1022] =  12'b000110101100; // 428
storage[1023] = -12'b000000010110; // -22
storage[1024] =  12'b000011101011; // 235
storage[1025] =  12'b000100011101; // 285
storage[1026] = -12'b000010101110; // -174
storage[1027] = -12'b000000101111; // -47
storage[1028] = -12'b000101011011; // -347
storage[1029] =  12'b000110110100; // 436
storage[1030] = -12'b000010111010; // -186
storage[1031] = -12'b000010110110; // -182
storage[1032] =  12'b000010011100; // 156
storage[1033] =  12'b000100011101; // 285
storage[1034] =  12'b001001000101; // 581
storage[1035] =  12'b000110101101; // 429
storage[1036] =  12'b001101100100; // 868
storage[1037] =  12'b001001101010; // 618
storage[1038] =  12'b000000010111; // 23
storage[1039] = -12'b000100110110; // -310
storage[1040] = -12'b001010011010; // -666
storage[1041] = -12'b000111010111; // -471
storage[1042] = -12'b000010110110; // -182
storage[1043] = -12'b000000001101; // -13
storage[1044] = -12'b000000011101; // -29
storage[1045] =  12'b000011001000; // 200
storage[1046] =  12'b000100111110; // 318
storage[1047] =  12'b001001100100; // 612
storage[1048] =  12'b000001100001; // 97
storage[1049] =  12'b000001111101; // 125
storage[1050] =  12'b000111111111; // 511
storage[1051] = -12'b001100111110; // -830
storage[1052] = -12'b000010100111; // -167
storage[1053] =  12'b000010000111; // 135
storage[1054] = -12'b000110010001; // -401
storage[1055] = -12'b000101100010; // -354
storage[1056] =  12'b000001000111; // 71
storage[1057] =  12'b000100110010; // 306
storage[1058] = -12'b000001000100; // -68
storage[1059] =  12'b000001100100; // 100
storage[1060] =  12'b000100000010; // 258
storage[1061] = -12'b000010001010; // -138
storage[1062] =  12'b000000001000; // 8
storage[1063] = -12'b000011000111; // -199
storage[1064] = -12'b000010100000; // -160
storage[1065] =  12'b000001100111; // 103
storage[1066] =  12'b000001011010; // 90
storage[1067] = -12'b001000010001; // -529
storage[1068] =  12'b000011001010; // 202
storage[1069] =  12'b000111011101; // 477
storage[1070] =  12'b000101011001; // 345
storage[1071] =  12'b000011011101; // 221
storage[1072] = -12'b001101110001; // -881
storage[1073] = -12'b000011011000; // -216
storage[1074] =  12'b000011100011; // 227
storage[1075] =  12'b000001111000; // 120
storage[1076] = -12'b000001101000; // -104
storage[1077] = -12'b000001110000; // -112
storage[1078] =  12'b000110101101; // 429
storage[1079] =  12'b000001000101; // 69
storage[1080] = -12'b000010110010; // -178
storage[1081] = -12'b000010000011; // -131
storage[1082] = -12'b001001001110; // -590
storage[1083] = -12'b000111100110; // -486
storage[1084] =  12'b000111010011; // 467
storage[1085] = -12'b000011000011; // -195
storage[1086] = -12'b010000100100; // -1060
storage[1087] =  12'b001010110110; // 694
storage[1088] =  12'b001011011001; // 729
storage[1089] =  12'b000100001010; // 266
storage[1090] =  12'b000110011000; // 408
storage[1091] =  12'b000100101011; // 299
storage[1092] =  12'b001001010010; // 594
storage[1093] = -12'b000110110100; // -436
storage[1094] = -12'b000101011100; // -348
storage[1095] =  12'b000010110011; // 179
storage[1096] = -12'b000101100000; // -352
storage[1097] = -12'b000101101010; // -362
storage[1098] = -12'b000110011000; // -408
storage[1099] =  12'b000101001000; // 328
storage[1100] =  12'b000011111001; // 249
storage[1101] = -12'b000000111010; // -58
storage[1102] =  12'b000111011011; // 475
storage[1103] =  12'b001010000100; // 644
storage[1104] =  12'b000001010101; // 85
storage[1105] = -12'b001000011011; // -539
storage[1106] =  12'b000001001000; // 72
storage[1107] =  12'b000101000111; // 327
storage[1108] =  12'b000001000100; // 68
storage[1109] = -12'b000000000011; // -3
storage[1110] = -12'b000000100110; // -38
storage[1111] = -12'b000010000101; // -133
storage[1112] = -12'b000010011000; // -152
storage[1113] =  12'b000100001110; // 270
storage[1114] = -12'b000011101000; // -232
storage[1115] = -12'b000001001111; // -79
storage[1116] =  12'b000101100100; // 356
storage[1117] = -12'b000000111000; // -56
storage[1118] =  12'b000000110101; // 53
storage[1119] =  12'b000010101100; // 172
storage[1120] =  12'b000100011100; // 284
storage[1121] =  12'b001001001100; // 588
storage[1122] =  12'b001100111110; // 830
storage[1123] =  12'b000101100000; // 352
storage[1124] =  12'b010000100001; // 1057
storage[1125] =  12'b001001101110; // 622
storage[1126] = -12'b000011100001; // -225
storage[1127] = -12'b000001111101; // -125
storage[1128] =  12'b000000000110; // 6
storage[1129] =  12'b000000101101; // 45
storage[1130] = -12'b000110001110; // -398
storage[1131] = -12'b000011010000; // -208
storage[1132] =  12'b000111101110; // 494
storage[1133] =  12'b000010000001; // 129
storage[1134] =  12'b000001000011; // 67
storage[1135] =  12'b000001100000; // 96
storage[1136] =  12'b000001110101; // 117
storage[1137] =  12'b000001011110; // 94
storage[1138] =  12'b000001001100; // 76
storage[1139] =  12'b000010100100; // 164
storage[1140] =  12'b000001000111; // 71
storage[1141] = -12'b001011000010; // -706
storage[1142] = -12'b001000001010; // -522
storage[1143] =  12'b000011011110; // 222
storage[1144] =  12'b000111000011; // 451
storage[1145] =  12'b000001100010; // 98
storage[1146] =  12'b000011100100; // 228
storage[1147] = -12'b000110010101; // -405
storage[1148] = -12'b000101010010; // -338
storage[1149] = -12'b000010101100; // -172
storage[1150] = -12'b010000100101; // -1061
storage[1151] = -12'b001111111111; // -1023
storage[1152] = -12'b000101100011; // -355
storage[1153] =  12'b000011011111; // 223
storage[1154] =  12'b000011001101; // 205
storage[1155] = -12'b000001111001; // -121
storage[1156] = -12'b000000101111; // -47
storage[1157] =  12'b000001100110; // 102
storage[1158] =  12'b000010001000; // 136
storage[1159] = -12'b000100101101; // -301
storage[1160] =  12'b000101010111; // 343
storage[1161] =  12'b001000001100; // 524
storage[1162] = -12'b000010111000; // -184
storage[1163] =  12'b000000000110; // 6
storage[1164] =  12'b000000000100; // 4
storage[1165] =  12'b000100100101; // 293
storage[1166] =  12'b000001110010; // 114
storage[1167] =  12'b000001111100; // 124
storage[1168] =  12'b000010011111; // 159
storage[1169] =  12'b000001001101; // 77
storage[1170] =  12'b000010011111; // 159
storage[1171] =  12'b000110000000; // 384
storage[1172] =  12'b000011110100; // 244
storage[1173] =  12'b000001001010; // 74
storage[1174] = -12'b000001011111; // -95
storage[1175] = -12'b001101100011; // -867
storage[1176] = -12'b001111000110; // -966
storage[1177] =  12'b000110010101; // 405
storage[1178] = -12'b000010110001; // -177
storage[1179] = -12'b010011100100; // -1252
storage[1180] =  12'b000111000100; // 452
storage[1181] =  12'b000001100110; // 102
storage[1182] =  12'b000001101100; // 108
storage[1183] =  12'b001100011010; // 794
storage[1184] =  12'b001010000101; // 645
storage[1185] =  12'b000110100100; // 420
storage[1186] =  12'b000101001011; // 331
storage[1187] =  12'b000001001101; // 77
storage[1188] =  12'b000001111100; // 124
storage[1189] = -12'b000000000101; // -5
storage[1190] =  12'b000010000100; // 132
storage[1191] = -12'b000111101111; // -495
storage[1192] = -12'b000010010100; // -148
storage[1193] = -12'b000101011110; // -350
storage[1194] =  12'b000000000011; // 3
storage[1195] = -12'b000000111101; // -61
storage[1196] =  12'b000001111000; // 120
storage[1197] =  12'b000001111111; // 127
storage[1198] =  12'b000100000011; // 259
storage[1199] =  12'b000011110011; // 243
storage[1200] =  12'b000010011011; // 155
storage[1201] =  12'b000000101011; // 43
storage[1202] = -12'b000001100010; // -98
storage[1203] = -12'b000101110111; // -375
storage[1204] =  12'b000010101101; // 173
storage[1205] = -12'b000100110110; // -310
storage[1206] =  12'b000011110100; // 244
storage[1207] = -12'b000100101110; // -302
storage[1208] =  12'b000110000110; // 390
storage[1209] =  12'b000011100101; // 229
storage[1210] = -12'b000000100101; // -37
storage[1211] =  12'b000000000100; // 4
storage[1212] =  12'b000010011010; // 154
storage[1213] =  12'b000010110001; // 177
storage[1214] =  12'b000001011100; // 92
storage[1215] =  12'b000100101000; // 296
storage[1216] = -12'b001001100001; // -609
storage[1217] = -12'b001000000001; // -513
storage[1218] =  12'b000110011011; // 411
storage[1219] = -12'b001001001100; // -588
storage[1220] =  12'b000000010001; // 17
storage[1221] =  12'b000101011010; // 346
storage[1222] =  12'b000001100010; // 98
storage[1223] =  12'b000010110110; // 182
storage[1224] = -12'b000000000110; // -6
storage[1225] =  12'b000100100110; // 294
storage[1226] =  12'b001000101110; // 558
storage[1227] = -12'b000001010111; // -87
storage[1228] =  12'b000001111110; // 126
storage[1229] =  12'b000111110110; // 502
storage[1230] =  12'b000100110100; // 308
storage[1231] =  12'b000010111010; // 186
storage[1232] =  12'b000011100110; // 230
storage[1233] =  12'b000001000010; // 66
storage[1234] =  12'b000001100111; // 103
storage[1235] =  12'b000001010010; // 82
storage[1236] =  12'b000010111101; // 189
storage[1237] =  12'b000001001011; // 75
storage[1238] = -12'b000101011001; // -345
storage[1239] = -12'b000000101001; // -41
storage[1240] = -12'b000100010010; // -274
storage[1241] = -12'b000011010101; // -213
storage[1242] =  12'b000011000000; // 192
storage[1243] =  12'b000110100000; // 416
storage[1244] =  12'b000110100101; // 421
storage[1245] = -12'b000000011100; // -28
storage[1246] =  12'b000010101111; // 175
storage[1247] =  12'b001011110111; // 759
storage[1248] =  12'b000111011000; // 472
storage[1249] =  12'b001011000001; // 705
storage[1250] =  12'b001100100110; // 806
storage[1251] =  12'b000011011100; // 220
storage[1252] = -12'b000010001111; // -143
storage[1253] =  12'b000010100101; // 165
storage[1254] =  12'b000100010110; // 278
storage[1255] = -12'b000011111000; // -248
storage[1256] = -12'b000010010011; // -147
storage[1257] =  12'b000010101010; // 170
storage[1258] = -12'b000101011011; // -347
storage[1259] = -12'b000001110001; // -113
storage[1260] =  12'b000000110110; // 54
storage[1261] = -12'b000100100010; // -290
storage[1262] = -12'b000000010111; // -23
storage[1263] =  12'b000101100000; // 352
storage[1264] =  12'b000000101010; // 42
storage[1265] = -12'b000000000100; // -4
storage[1266] = -12'b000001110111; // -119
storage[1267] =  12'b000100010001; // 273
storage[1268] =  12'b000011101101; // 237
storage[1269] = -12'b000000100101; // -37
storage[1270] =  12'b000111101101; // 493
storage[1271] =  12'b000100010011; // 275
storage[1272] =  12'b000100110000; // 304
storage[1273] =  12'b000100101100; // 300
storage[1274] =  12'b000111111100; // 508
storage[1275] =  12'b000101001000; // 328
storage[1276] =  12'b000100010111; // 279
storage[1277] =  12'b000100100100; // 292
storage[1278] = -12'b000000101001; // -41
storage[1279] =  12'b000000010010; // 18
storage[1280] = -12'b000011001010; // -202
storage[1281] =  12'b000010100001; // 161
storage[1282] = -12'b000001011101; // -93
storage[1283] =  12'b000001000101; // 69
storage[1284] =  12'b000000010001; // 17
storage[1285] =  12'b000000100101; // 37
storage[1286] = -12'b000101011011; // -347
storage[1287] =  12'b000000010000; // 16
storage[1288] = -12'b000010110001; // -177
storage[1289] = -12'b000010010101; // -149
storage[1290] =  12'b001000111111; // 575
storage[1291] =  12'b000001101010; // 106
storage[1292] = -12'b000001010100; // -84
storage[1293] =  12'b000001011010; // 90
storage[1294] =  12'b000010101101; // 173
storage[1295] =  12'b000001101010; // 106
storage[1296] = -12'b000010110011; // -179
storage[1297] = -12'b000110000011; // -387
storage[1298] =  12'b000000000000; // 0
storage[1299] =  12'b000010010111; // 151
storage[1300] = -12'b000110010010; // -402
storage[1301] = -12'b000001110110; // -118
storage[1302] = -12'b000000001100; // -12
storage[1303] = -12'b000100101000; // -296
storage[1304] = -12'b000011100100; // -228
storage[1305] =  12'b000011011100; // 220
storage[1306] =  12'b000010111010; // 186
storage[1307] = -12'b000000011111; // -31
storage[1308] = -12'b000001010110; // -86
storage[1309] =  12'b000011001011; // 203
storage[1310] =  12'b000000001001; // 9
storage[1311] = -12'b000010000111; // -135
storage[1312] = -12'b000001101010; // -106
storage[1313] = -12'b000000100110; // -38
storage[1314] =  12'b000000010100; // 20
storage[1315] =  12'b000011101110; // 238
storage[1316] =  12'b000010110000; // 176
storage[1317] =  12'b000001110010; // 114
storage[1318] =  12'b000100000011; // 259
storage[1319] =  12'b000101111001; // 377
storage[1320] =  12'b000110010010; // 402
storage[1321] =  12'b000000111111; // 63
storage[1322] =  12'b000000111011; // 59
storage[1323] =  12'b000000011001; // 25
storage[1324] = -12'b000001000100; // -68
storage[1325] = -12'b000011000100; // -196
storage[1326] = -12'b000010101101; // -173
storage[1327] = -12'b000011011010; // -218
storage[1328] = -12'b001000010111; // -535
storage[1329] = -12'b001011010101; // -725
storage[1330] = -12'b000000010100; // -20
storage[1331] =  12'b000100000011; // 259
storage[1332] =  12'b000001011010; // 90
storage[1333] =  12'b000011001011; // 203
storage[1334] = -12'b000100001001; // -265
storage[1335] = -12'b000100101110; // -302
storage[1336] = -12'b000000110110; // -54
storage[1337] =  12'b000100000111; // 263
storage[1338] = -12'b000000110010; // -50
storage[1339] =  12'b000010010110; // 150
storage[1340] =  12'b000100000100; // 260
storage[1341] =  12'b000100010001; // 273
storage[1342] =  12'b000100001011; // 267
storage[1343] =  12'b000010011101; // 157
storage[1344] = -12'b000000000101; // -5
storage[1345] =  12'b000000100001; // 33
storage[1346] =  12'b000101000010; // 322
storage[1347] = -12'b000000101010; // -42
storage[1348] = -12'b000010101101; // -173
storage[1349] =  12'b000010010001; // 145
storage[1350] =  12'b000101001111; // 335
storage[1351] =  12'b000000011010; // 26
storage[1352] =  12'b000110111110; // 446
storage[1353] =  12'b001011010110; // 726
storage[1354] = -12'b000010000000; // -128
storage[1355] =  12'b000011111010; // 250
storage[1356] =  12'b001100110101; // 821
storage[1357] =  12'b000111000101; // 453
storage[1358] = -12'b000110100111; // -423
storage[1359] = -12'b000011110110; // -246
storage[1360] =  12'b000011001101; // 205
storage[1361] =  12'b000110101101; // 429
storage[1362] =  12'b001000101110; // 558
storage[1363] = -12'b000001000001; // -65
storage[1364] =  12'b000000110011; // 51
storage[1365] =  12'b001011001010; // 714
storage[1366] = -12'b000000001001; // -9
storage[1367] = -12'b000100010010; // -274
storage[1368] =  12'b000110101010; // 426
storage[1369] =  12'b000001100110; // 102
storage[1370] =  12'b000001011111; // 95
storage[1371] = -12'b000001001111; // -79
storage[1372] = -12'b000011111111; // -255
storage[1373] =  12'b000100100011; // 291
storage[1374] = -12'b000000100101; // -37
storage[1375] = -12'b000011000001; // -193
storage[1376] = -12'b000010101001; // -169
storage[1377] = -12'b000011100001; // -225
storage[1378] =  12'b000100100111; // 295
storage[1379] =  12'b000001010100; // 84
storage[1380] = -12'b000001101111; // -111
storage[1381] = -12'b000001010000; // -80
storage[1382] =  12'b000001101010; // 106
storage[1383] = -12'b000100001101; // -269
storage[1384] =  12'b000010011001; // 153
storage[1385] = -12'b000001111011; // -123
storage[1386] = -12'b000001011101; // -93
storage[1387] = -12'b000010011110; // -158
storage[1388] = -12'b000010111110; // -190
storage[1389] = -12'b000001101100; // -108
storage[1390] = -12'b000100010100; // -276
storage[1391] = -12'b000011111011; // -251
storage[1392] =  12'b000100111111; // 319
storage[1393] = -12'b000010100101; // -165
storage[1394] = -12'b000110100100; // -420
storage[1395] =  12'b000000001001; // 9
storage[1396] = -12'b000111100000; // -480
storage[1397] =  12'b000100100111; // 295
storage[1398] =  12'b001000000010; // 514
storage[1399] =  12'b000010001011; // 139
storage[1400] = -12'b000001100001; // -97
storage[1401] = -12'b000111100110; // -486
storage[1402] =  12'b000110100010; // 418
storage[1403] = -12'b000111011011; // -475
storage[1404] = -12'b001000110001; // -561
storage[1405] =  12'b000010001000; // 136
storage[1406] =  12'b000100000011; // 259
storage[1407] = -12'b000000011100; // -28
storage[1408] =  12'b000011100011; // 227
storage[1409] =  12'b000001101100; // 108
storage[1410] = -12'b000110100001; // -417
storage[1411] =  12'b000010101110; // 174
storage[1412] = -12'b000010000001; // -129
storage[1413] = -12'b001000011000; // -536
storage[1414] = -12'b000010111011; // -187
storage[1415] =  12'b000111101100; // 492
storage[1416] = -12'b000100000100; // -260
storage[1417] =  12'b001000001111; // 527
storage[1418] =  12'b000111010110; // 470
storage[1419] = -12'b001010011100; // -668
storage[1420] =  12'b000101101111; // 367
storage[1421] = -12'b000001011000; // -88
storage[1422] = -12'b001000001101; // -525
storage[1423] =  12'b000110100001; // 417
storage[1424] = -12'b000000001101; // -13
storage[1425] = -12'b000010011110; // -158
storage[1426] = -12'b000110011110; // -414
storage[1427] = -12'b000110101100; // -428
storage[1428] = -12'b001000101001; // -553
storage[1429] = -12'b000100111000; // -312
storage[1430] = -12'b000001111100; // -124
storage[1431] = -12'b000110000010; // -386
storage[1432] = -12'b000100001100; // -268
storage[1433] =  12'b000100111001; // 313
storage[1434] =  12'b000001011100; // 92
storage[1435] =  12'b000011110110; // 246
storage[1436] =  12'b000101000000; // 320
storage[1437] = -12'b001011000101; // -709
storage[1438] =  12'b000111010010; // 466
storage[1439] = -12'b000000011001; // -25
storage[1440] = -12'b001000001101; // -525
storage[1441] = -12'b000000011100; // -28
storage[1442] =  12'b000010100111; // 167
storage[1443] = -12'b000010100101; // -165
storage[1444] =  12'b000000011011; // 27
storage[1445] = -12'b001011010110; // -726
storage[1446] = -12'b001001100000; // -608
storage[1447] = -12'b000011010111; // -215
storage[1448] = -12'b010000110010; // -1074
storage[1449] =  12'b000111001101; // 461
storage[1450] = -12'b000000101100; // -44
storage[1451] =  12'b000100110000; // 304
storage[1452] = -12'b000010111101; // -189
storage[1453] = -12'b000100101001; // -297
storage[1454] =  12'b000100011010; // 282
storage[1455] =  12'b000111001100; // 460
storage[1456] =  12'b000000110011; // 51
storage[1457] =  12'b000110001001; // 393
storage[1458] = -12'b000001110001; // -113
storage[1459] = -12'b000100001000; // -264
storage[1460] = -12'b000110001111; // -399
storage[1461] =  12'b000010110001; // 177
storage[1462] = -12'b001001001011; // -587
storage[1463] =  12'b000100110100; // 308
storage[1464] =  12'b000101011111; // 351
storage[1465] =  12'b000010101110; // 174
storage[1466] =  12'b000110111101; // 445
storage[1467] = -12'b000010001110; // -142
storage[1468] =  12'b000110000011; // 387
storage[1469] = -12'b000000011010; // -26
storage[1470] = -12'b000011011011; // -219
storage[1471] =  12'b001010110010; // 690
storage[1472] = -12'b000001010101; // -85
storage[1473] = -12'b000100011101; // -285
storage[1474] =  12'b010001111011; // 1147
storage[1475] = -12'b000101100111; // -359
storage[1476] = -12'b000101011110; // -350
storage[1477] =  12'b000011101001; // 233
storage[1478] = -12'b001011011001; // -729
storage[1479] = -12'b000110100111; // -423
storage[1480] =  12'b000001010000; // 80
storage[1481] = -12'b001011100110; // -742
storage[1482] = -12'b000011111110; // -254
storage[1483] =  12'b000101010100; // 340
storage[1484] = -12'b000110110100; // -436
storage[1485] =  12'b000001000100; // 68
storage[1486] = -12'b000001110101; // -117
storage[1487] = -12'b000100111000; // -312
storage[1488] = -12'b000000010001; // -17
storage[1489] =  12'b000001100010; // 98
storage[1490] = -12'b000100101111; // -303
storage[1491] =  12'b000010101100; // 172
storage[1492] =  12'b000010011110; // 158
storage[1493] = -12'b000100100011; // -291
storage[1494] = -12'b000001111101; // -125
storage[1495] =  12'b000010010001; // 145
storage[1496] = -12'b000011001110; // -206
storage[1497] = -12'b000100101010; // -298
storage[1498] = -12'b000001110010; // -114
storage[1499] = -12'b000001100011; // -99
storage[1500] = -12'b000110001001; // -393
storage[1501] =  12'b000000111000; // 56
storage[1502] = -12'b000001111000; // -120
storage[1503] = -12'b000000001111; // -15
storage[1504] =  12'b000100001011; // 267
storage[1505] = -12'b000100100000; // -288
storage[1506] = -12'b000101001010; // -330
storage[1507] =  12'b000000110001; // 49
storage[1508] = -12'b000101000001; // -321
storage[1509] = -12'b000011001010; // -202
storage[1510] = -12'b000000001000; // -8
storage[1511] =  12'b000100100111; // 295
storage[1512] =  12'b000000001001; // 9
storage[1513] =  12'b000010100000; // 160
storage[1514] = -12'b000010010110; // -150
storage[1515] = -12'b000011010000; // -208
storage[1516] = -12'b000010110000; // -176
storage[1517] = -12'b000000010101; // -21
storage[1518] = -12'b000000100110; // -38
storage[1519] = -12'b000010011001; // -153
storage[1520] = -12'b000001111010; // -122
storage[1521] = -12'b000000100000; // -32
storage[1522] =  12'b000000101101; // 45
storage[1523] =  12'b000001111000; // 120
storage[1524] =  12'b000010000111; // 135
storage[1525] = -12'b000000010111; // -23
storage[1526] =  12'b000001010110; // 86
storage[1527] =  12'b000010001100; // 140
storage[1528] = -12'b000000011101; // -29
storage[1529] = -12'b000010001101; // -141
storage[1530] =  12'b000100100001; // 289
storage[1531] =  12'b000101010110; // 342
storage[1532] =  12'b000010010100; // 148
storage[1533] =  12'b000011011010; // 218
storage[1534] =  12'b001001100111; // 615
storage[1535] =  12'b000111001100; // 460
storage[1536] =  12'b000001001001; // 73
storage[1537] =  12'b001001001001; // 585
storage[1538] =  12'b000011111010; // 250
storage[1539] =  12'b000110011010; // 410
storage[1540] =  12'b000100100111; // 295
storage[1541] = -12'b000010100101; // -165
storage[1542] =  12'b000000000101; // 5
storage[1543] =  12'b001011000010; // 706
storage[1544] =  12'b000010111101; // 189
storage[1545] = -12'b000001100110; // -102
storage[1546] = -12'b000001110010; // -114
storage[1547] = -12'b000001010101; // -85
storage[1548] =  12'b000001000001; // 65
storage[1549] =  12'b000001101101; // 109
storage[1550] = -12'b000010100110; // -166
storage[1551] = -12'b000000010010; // -18
storage[1552] = -12'b000001100001; // -97
storage[1553] = -12'b000001010100; // -84
storage[1554] = -12'b000011001001; // -201
storage[1555] = -12'b000111011100; // -476
storage[1556] = -12'b001101100100; // -868
storage[1557] = -12'b000011100010; // -226
storage[1558] =  12'b000000101001; // 41
storage[1559] =  12'b000011100110; // 230
storage[1560] = -12'b000011110110; // -246
storage[1561] =  12'b000100111010; // 314
storage[1562] = -12'b000100000110; // -262
storage[1563] = -12'b000000000110; // -6
storage[1564] = -12'b001000101001; // -553
storage[1565] = -12'b001001110110; // -630
storage[1566] =  12'b000101110001; // 369
storage[1567] =  12'b000101001100; // 332
storage[1568] =  12'b000110110011; // 435
storage[1569] =  12'b001010011010; // 666
storage[1570] = -12'b000111110101; // -501
storage[1571] = -12'b000100110110; // -310
storage[1572] =  12'b000000001110; // 14
storage[1573] =  12'b000001010010; // 82
storage[1574] =  12'b000010010101; // 149
storage[1575] =  12'b000111101101; // 493
storage[1576] = -12'b000011011100; // -220
storage[1577] = -12'b000001000000; // -64
storage[1578] = -12'b000000101000; // -40
storage[1579] = -12'b001010000101; // -645
storage[1580] = -12'b001001001100; // -588
storage[1581] = -12'b000100100010; // -290
storage[1582] = -12'b001010000110; // -646
storage[1583] = -12'b000111011011; // -475
storage[1584] = -12'b000001101100; // -108
storage[1585] =  12'b000000010010; // 18
storage[1586] =  12'b000100010010; // 274
storage[1587] = -12'b000100000001; // -257
storage[1588] = -12'b000010011110; // -158
storage[1589] = -12'b000011101111; // -239
storage[1590] = -12'b000110000110; // -390
storage[1591] = -12'b001010111011; // -699
storage[1592] = -12'b001001100010; // -610
storage[1593] = -12'b000001001110; // -78
storage[1594] =  12'b000100100101; // 293
storage[1595] = -12'b000001010101; // -85
storage[1596] = -12'b000001100011; // -99
storage[1597] =  12'b000001101001; // 105
storage[1598] =  12'b000100110110; // 310
storage[1599] =  12'b000101011011; // 347
storage[1600] =  12'b000100001010; // 266
storage[1601] =  12'b000100000010; // 258
storage[1602] =  12'b000110110111; // 439
storage[1603] =  12'b000000011000; // 24
storage[1604] = -12'b000000001111; // -15
storage[1605] =  12'b000011010110; // 214
storage[1606] =  12'b000000100001; // 33
storage[1607] =  12'b000000111111; // 63
storage[1608] =  12'b000101001111; // 335
storage[1609] =  12'b000110111110; // 446
storage[1610] =  12'b000010001101; // 141
storage[1611] =  12'b000001011000; // 88
storage[1612] = -12'b000010110001; // -177
storage[1613] = -12'b000110010100; // -404
storage[1614] =  12'b000000100001; // 33
storage[1615] = -12'b000000011010; // -26
storage[1616] =  12'b000011100100; // 228
storage[1617] =  12'b000011101111; // 239
storage[1618] =  12'b000010010111; // 151
storage[1619] =  12'b000001101101; // 109
storage[1620] =  12'b000001010011; // 83
storage[1621] = -12'b000111000010; // -450
storage[1622] = -12'b000001001001; // -73
storage[1623] =  12'b000000010101; // 21
storage[1624] =  12'b000100011000; // 280
storage[1625] =  12'b000001111001; // 121
storage[1626] =  12'b000011111011; // 251
storage[1627] = -12'b000010010101; // -149
storage[1628] = -12'b000010001010; // -138
storage[1629] = -12'b000100110111; // -311
storage[1630] =  12'b001001001010; // 586
storage[1631] =  12'b001001110010; // 626
storage[1632] =  12'b000110010011; // 403
storage[1633] =  12'b001001111110; // 638
storage[1634] =  12'b001100101101; // 813
storage[1635] =  12'b000000011001; // 25
storage[1636] = -12'b000011010101; // -213
storage[1637] = -12'b000001010110; // -86
storage[1638] = -12'b000101010101; // -341
storage[1639] = -12'b000001101011; // -107
storage[1640] =  12'b000000000100; // 4
storage[1641] =  12'b000011011011; // 219
storage[1642] = -12'b000100010101; // -277
storage[1643] = -12'b001001101111; // -623
storage[1644] = -12'b000001010111; // -87
storage[1645] =  12'b000010011011; // 155
storage[1646] =  12'b000110011010; // 410
storage[1647] =  12'b001000010111; // 535
storage[1648] = -12'b000011001111; // -207
storage[1649] = -12'b000000001010; // -10
storage[1650] = -12'b001000001101; // -525
storage[1651] =  12'b000101101000; // 360
storage[1652] = -12'b000000010111; // -23
storage[1653] =  12'b000001101110; // 110
storage[1654] =  12'b000001010101; // 85
storage[1655] = -12'b000100111010; // -314
storage[1656] = -12'b000011011101; // -221
storage[1657] = -12'b000111101010; // -490
storage[1658] =  12'b000001010001; // 81
storage[1659] =  12'b000001000000; // 64
storage[1660] =  12'b000010110001; // 177
storage[1661] = -12'b000001110011; // -115
storage[1662] =  12'b000001100101; // 101
storage[1663] = -12'b000000011101; // -29
storage[1664] =  12'b000011011100; // 220
storage[1665] = -12'b000000001010; // -10
storage[1666] =  12'b000000001110; // 14
storage[1667] =  12'b000110001111; // 399
storage[1668] = -12'b000010110011; // -179
storage[1669] =  12'b000001100000; // 96
storage[1670] = -12'b000000110011; // -51
storage[1671] =  12'b000100110111; // 311
storage[1672] =  12'b000110111010; // 442
storage[1673] = -12'b000001001111; // -79
storage[1674] =  12'b000100001110; // 270
storage[1675] =  12'b000001101101; // 109
storage[1676] = -12'b000111011001; // -473
storage[1677] = -12'b000101110001; // -369
storage[1678] = -12'b000100101111; // -303
storage[1679] = -12'b000011110011; // -243
storage[1680] =  12'b000000101101; // 45
storage[1681] =  12'b000010110100; // 180
storage[1682] =  12'b000001001010; // 74
storage[1683] = -12'b000000101101; // -45
storage[1684] =  12'b000101010001; // 337
storage[1685] = -12'b000001001110; // -78
storage[1686] = -12'b000010001100; // -140
storage[1687] =  12'b000011001010; // 202
storage[1688] =  12'b000001111100; // 124
storage[1689] =  12'b000101110000; // 368
storage[1690] =  12'b000011100010; // 226
storage[1691] =  12'b000100011101; // 285
storage[1692] =  12'b000101011011; // 347
storage[1693] =  12'b000011011101; // 221
storage[1694] =  12'b000011111001; // 249
storage[1695] =  12'b000010100110; // 166
storage[1696] =  12'b000000010110; // 22
storage[1697] =  12'b000011000001; // 193
storage[1698] =  12'b000110001010; // 394
storage[1699] =  12'b000100011111; // 287
storage[1700] =  12'b000011110011; // 243
storage[1701] =  12'b001010101011; // 683
storage[1702] = -12'b000101011100; // -348
storage[1703] = -12'b000010001001; // -137
storage[1704] =  12'b000010100110; // 166
storage[1705] = -12'b000001001001; // -73
storage[1706] = -12'b000111001001; // -457
storage[1707] =  12'b000010111011; // 187
storage[1708] =  12'b000001111010; // 122
storage[1709] = -12'b000000000110; // -6
storage[1710] = -12'b000000001111; // -15
storage[1711] = -12'b000100001011; // -267
storage[1712] = -12'b000111011000; // -472
storage[1713] = -12'b000000110100; // -52
storage[1714] = -12'b000110100110; // -422
storage[1715] = -12'b000111001000; // -456
storage[1716] = -12'b001010001111; // -655
storage[1717] = -12'b000110100001; // -417
storage[1718] =  12'b000010011111; // 159
storage[1719] = -12'b000011110000; // -240
storage[1720] = -12'b000010001110; // -142
storage[1721] = -12'b000111011100; // -476
storage[1722] = -12'b000100101010; // -298
storage[1723] = -12'b000011001101; // -205
storage[1724] = -12'b000110100101; // -421
storage[1725] = -12'b000000010111; // -23
storage[1726] =  12'b000100111101; // 317
storage[1727] =  12'b000011110100; // 244
storage[1728] =  12'b000100101111; // 303
storage[1729] = -12'b000100011010; // -282
storage[1730] = -12'b000000000110; // -6
storage[1731] = -12'b000010111101; // -189
storage[1732] =  12'b000001000001; // 65
storage[1733] =  12'b000001000010; // 66
storage[1734] =  12'b000010100101; // 165
storage[1735] = -12'b000100000001; // -257
storage[1736] =  12'b000100001100; // 268
storage[1737] =  12'b001001000101; // 581
storage[1738] = -12'b000110010100; // -404
storage[1739] = -12'b000000011111; // -31
storage[1740] = -12'b000000101101; // -45
storage[1741] = -12'b000000000100; // -4
storage[1742] = -12'b000011111110; // -254
storage[1743] =  12'b000000000111; // 7
storage[1744] =  12'b000001101110; // 110
storage[1745] =  12'b000110001110; // 398
storage[1746] =  12'b000101101100; // 364
storage[1747] = -12'b000001111001; // -121
storage[1748] = -12'b000010111111; // -191
storage[1749] = -12'b000011111101; // -253
storage[1750] = -12'b000011010100; // -212
storage[1751] =  12'b000001100101; // 101
storage[1752] = -12'b000001101111; // -111
storage[1753] =  12'b000100000111; // 263
storage[1754] =  12'b000011100010; // 226
storage[1755] =  12'b000000100011; // 35
storage[1756] =  12'b000000011011; // 27
storage[1757] =  12'b000101010101; // 341
storage[1758] =  12'b000010110110; // 182
storage[1759] = -12'b000101100100; // -356
storage[1760] =  12'b000100001000; // 264
storage[1761] = -12'b000000101111; // -47
storage[1762] = -12'b000000111111; // -63
storage[1763] = -12'b000001100011; // -99
storage[1764] = -12'b000001100110; // -102
storage[1765] = -12'b000001101001; // -105
storage[1766] =  12'b000000100110; // 38
storage[1767] =  12'b000011110101; // 245
storage[1768] = -12'b000000011111; // -31
storage[1769] =  12'b000001000110; // 70
storage[1770] =  12'b000010010101; // 149
storage[1771] = -12'b000011001001; // -201
storage[1772] =  12'b000001101101; // 109
storage[1773] =  12'b000001000100; // 68
storage[1774] = -12'b000001111111; // -127
storage[1775] = -12'b000000110010; // -50
storage[1776] =  12'b000000010101; // 21
storage[1777] = -12'b000001011110; // -94
storage[1778] =  12'b000001101011; // 107
storage[1779] = -12'b000011001110; // -206
storage[1780] = -12'b000100001010; // -266
storage[1781] = -12'b000000111011; // -59
storage[1782] = -12'b000001101100; // -108
storage[1783] =  12'b001000000111; // 519
storage[1784] = -12'b001101010111; // -855
storage[1785] = -12'b001100010001; // -785
storage[1786] = -12'b001000001100; // -524
storage[1787] = -12'b011101000110; // -1862
storage[1788] = -12'b000010001111; // -143
storage[1789] = -12'b010101111000; // -1400
storage[1790] = -12'b001000001011; // -523
storage[1791] =  12'b000111001111; // 463
storage[1792] =  12'b000110010000; // 400
storage[1793] = -12'b000100101100; // -300
storage[1794] = -12'b000010110101; // -181
storage[1795] = -12'b000011011100; // -220
storage[1796] = -12'b000001011010; // -90
storage[1797] =  12'b000010011101; // 157
storage[1798] =  12'b000111011111; // 479
storage[1799] =  12'b000000101110; // 46
storage[1800] =  12'b000111001011; // 459
storage[1801] =  12'b000010101101; // 173
storage[1802] =  12'b000101000000; // 320
storage[1803] =  12'b000110101011; // 427
storage[1804] =  12'b000010001110; // 142
storage[1805] =  12'b000101100100; // 356
storage[1806] = -12'b000001111000; // -120
storage[1807] = -12'b000010001100; // -140
storage[1808] =  12'b000000110111; // 55
storage[1809] =  12'b000010100000; // 160
storage[1810] =  12'b000110010100; // 404
storage[1811] =  12'b000010011100; // 156
storage[1812] = -12'b000010011000; // -152
storage[1813] = -12'b000001110111; // -119
storage[1814] =  12'b000101001010; // 330
storage[1815] = -12'b000000110101; // -53
storage[1816] =  12'b000000010011; // 19
storage[1817] = -12'b000100111001; // -313
storage[1818] =  12'b000011100101; // 229
storage[1819] =  12'b001000001110; // 526
storage[1820] =  12'b000000001000; // 8
storage[1821] = -12'b000001111101; // -125
storage[1822] = -12'b000011111101; // -253
storage[1823] =  12'b000001101111; // 111
storage[1824] =  12'b000001101100; // 108
storage[1825] = -12'b001001101110; // -622
storage[1826] =  12'b000100100100; // 292
storage[1827] =  12'b001010010011; // 659
storage[1828] =  12'b000011111110; // 254
storage[1829] =  12'b000001010010; // 82
storage[1830] = -12'b000001001011; // -75
storage[1831] = -12'b000100110001; // -305
storage[1832] = -12'b000010111111; // -191
storage[1833] = -12'b000100111001; // -313
storage[1834] =  12'b000001000010; // 66
storage[1835] =  12'b000100111011; // 315
storage[1836] =  12'b000110000110; // 390
storage[1837] =  12'b000101001010; // 330
storage[1838] = -12'b000001010111; // -87
storage[1839] = -12'b000110000101; // -389
storage[1840] = -12'b000001010111; // -87
storage[1841] = -12'b000101101001; // -361
storage[1842] = -12'b000110110000; // -432
storage[1843] =  12'b000100110011; // 307
storage[1844] =  12'b000011100101; // 229
storage[1845] =  12'b000001010100; // 84
storage[1846] = -12'b000010000100; // -132
storage[1847] = -12'b000010101101; // -173
storage[1848] =  12'b000001010111; // 87
storage[1849] = -12'b000101010011; // -339
storage[1850] = -12'b001011001001; // -713
storage[1851] = -12'b001101101001; // -873
storage[1852] = -12'b000010000000; // -128
storage[1853] = -12'b000011111111; // -255
storage[1854] = -12'b000111100110; // -486
storage[1855] =  12'b000101101110; // 366
storage[1856] = -12'b000000101110; // -46
storage[1857] = -12'b000001100011; // -99
storage[1858] = -12'b000010000101; // -133
storage[1859] =  12'b000001111100; // 124
storage[1860] = -12'b000101010011; // -339
storage[1861] =  12'b000011000110; // 198
storage[1862] =  12'b000011001101; // 205
storage[1863] = -12'b000000000100; // -4
storage[1864] =  12'b000000001111; // 15
storage[1865] =  12'b000010010110; // 150
storage[1866] =  12'b000000001111; // 15
storage[1867] =  12'b000110011010; // 410
storage[1868] =  12'b000010101111; // 175
storage[1869] = -12'b000000011101; // -29
storage[1870] =  12'b000110001100; // 396
storage[1871] =  12'b000010100001; // 161
storage[1872] =  12'b000000111011; // 59
storage[1873] =  12'b000010101110; // 174
storage[1874] = -12'b000011010011; // -211
storage[1875] = -12'b000010111101; // -189
storage[1876] =  12'b000011001010; // 202
storage[1877] =  12'b000010101110; // 174
storage[1878] =  12'b000001111011; // 123
storage[1879] =  12'b000000110101; // 53
storage[1880] = -12'b000010010100; // -148
storage[1881] =  12'b000001010011; // 83
storage[1882] =  12'b000010110101; // 181
storage[1883] =  12'b000000000011; // 3
storage[1884] = -12'b000100111101; // -317
storage[1885] =  12'b000010110110; // 182
storage[1886] =  12'b000010001011; // 139
storage[1887] =  12'b000010010010; // 146
storage[1888] = -12'b000010110000; // -176
storage[1889] =  12'b000001101110; // 110
storage[1890] =  12'b000100111110; // 318
storage[1891] =  12'b000100011010; // 282
storage[1892] = -12'b000000000010; // -2
storage[1893] =  12'b000000100100; // 36
storage[1894] =  12'b000010100111; // 167
storage[1895] =  12'b000011111100; // 252
storage[1896] = -12'b000001111000; // -120
storage[1897] =  12'b000000000001; // 1
storage[1898] = -12'b000011111101; // -253
storage[1899] = -12'b000011110010; // -242
storage[1900] = -12'b000100001001; // -265
storage[1901] = -12'b000010001011; // -139
storage[1902] = -12'b000010111001; // -185
storage[1903] = -12'b000010111111; // -191
storage[1904] = -12'b000101011111; // -351
storage[1905] = -12'b000001111100; // -124
storage[1906] =  12'b000000100101; // 37
storage[1907] = -12'b000010001100; // -140
storage[1908] = -12'b000010010110; // -150
storage[1909] = -12'b000001010110; // -86
storage[1910] =  12'b000010000001; // 129
storage[1911] =  12'b000001010010; // 82
storage[1912] = -12'b000000101100; // -44
storage[1913] =  12'b000001111010; // 122
storage[1914] = -12'b000000001000; // -8
storage[1915] =  12'b000011100100; // 228
storage[1916] =  12'b000010101001; // 169
storage[1917] =  12'b000010110011; // 179
storage[1918] = -12'b000011000100; // -196
storage[1919] = -12'b000000101101; // -45
storage[1920] =  12'b000101110110; // 374
storage[1921] = -12'b000010010111; // -151
storage[1922] = -12'b000000010011; // -19
storage[1923] = -12'b000000100100; // -36
storage[1924] =  12'b000011101111; // 239
storage[1925] =  12'b000011101111; // 239
storage[1926] =  12'b000000100011; // 35
storage[1927] = -12'b000100100100; // -292
storage[1928] = -12'b000001111011; // -123
storage[1929] =  12'b000110001011; // 395
storage[1930] = -12'b000101100110; // -358
storage[1931] = -12'b000100101111; // -303
storage[1932] =  12'b000010011101; // 157
storage[1933] =  12'b000100011100; // 284
storage[1934] =  12'b000001111101; // 125
storage[1935] =  12'b000100001001; // 265
storage[1936] = -12'b001001101001; // -617
storage[1937] = -12'b000011100011; // -227
storage[1938] =  12'b000010000011; // 131
storage[1939] = -12'b000010101101; // -173
storage[1940] = -12'b000001010000; // -80
storage[1941] =  12'b000001111111; // 127
storage[1942] =  12'b000001000010; // 66
storage[1943] =  12'b000011010110; // 214
storage[1944] =  12'b000100101011; // 299
storage[1945] = -12'b000011011110; // -222
storage[1946] =  12'b000011010110; // 214
storage[1947] =  12'b000110110110; // 438
storage[1948] =  12'b000001101101; // 109
storage[1949] =  12'b000010010101; // 149
storage[1950] =  12'b000100000110; // 262
storage[1951] =  12'b000010011001; // 153
storage[1952] =  12'b000010000000; // 128
storage[1953] =  12'b000000110111; // 55
storage[1954] =  12'b000010001110; // 142
storage[1955] =  12'b000001011100; // 92
storage[1956] = -12'b000011101110; // -238
storage[1957] =  12'b000001000000; // 64
storage[1958] = -12'b000000010101; // -21
storage[1959] =  12'b000000010011; // 19
storage[1960] = -12'b000000010111; // -23
storage[1961] = -12'b000010011001; // -153
storage[1962] = -12'b000000000001; // -1
storage[1963] =  12'b000001000001; // 65
storage[1964] =  12'b000001011000; // 88
storage[1965] =  12'b000010101000; // 168
storage[1966] =  12'b000000101011; // 43
storage[1967] =  12'b000010000100; // 132
storage[1968] = -12'b000010100011; // -163
storage[1969] =  12'b000000011110; // 30
storage[1970] = -12'b000001011101; // -93
storage[1971] = -12'b000010010000; // -144
storage[1972] =  12'b000011101101; // 237
storage[1973] =  12'b000011000011; // 195
storage[1974] =  12'b000010101001; // 169
storage[1975] =  12'b000000101011; // 43
storage[1976] = -12'b000000101100; // -44
storage[1977] = -12'b000101100111; // -359
storage[1978] =  12'b000010101010; // 170
storage[1979] =  12'b000010011110; // 158
storage[1980] =  12'b000000110110; // 54
storage[1981] = -12'b000001100101; // -101
storage[1982] =  12'b000001011101; // 93
storage[1983] =  12'b000010000010; // 130
storage[1984] = -12'b000001001011; // -75
storage[1985] =  12'b000010101111; // 175
storage[1986] = -12'b000011001100; // -204
storage[1987] =  12'b000010001101; // 141
storage[1988] =  12'b000001111110; // 126
storage[1989] = -12'b000100001010; // -266
storage[1990] =  12'b000001011111; // 95
storage[1991] =  12'b000001001010; // 74
storage[1992] =  12'b000010001001; // 137
storage[1993] = -12'b001000011100; // -540
storage[1994] = -12'b001100010110; // -790
storage[1995] = -12'b001101110111; // -887
storage[1996] = -12'b000001110100; // -116
storage[1997] = -12'b000100101110; // -302
storage[1998] = -12'b001010011000; // -664
storage[1999] =  12'b000011101010; // 234
storage[2000] =  12'b000010111110; // 190
storage[2001] =  12'b000001001001; // 73
storage[2002] =  12'b000001110010; // 114
storage[2003] = -12'b000101100111; // -359
storage[2004] = -12'b001000100111; // -551
storage[2005] = -12'b000000101101; // -45
storage[2006] = -12'b000010011011; // -155
storage[2007] = -12'b000000111110; // -62
storage[2008] =  12'b000011010111; // 215
storage[2009] =  12'b000010100011; // 163
storage[2010] =  12'b000001011001; // 89
storage[2011] = -12'b000001111101; // -125
storage[2012] = -12'b000010100000; // -160
storage[2013] = -12'b000100011000; // -280
storage[2014] = -12'b000100001001; // -265
storage[2015] = -12'b000011100110; // -230
storage[2016] = -12'b000011001101; // -205
storage[2017] = -12'b000000100010; // -34
storage[2018] =  12'b000001000110; // 70
storage[2019] =  12'b000001100000; // 96
storage[2020] =  12'b000011100110; // 230
storage[2021] =  12'b000010001011; // 139
storage[2022] =  12'b000100010011; // 275
storage[2023] =  12'b000000100001; // 33
storage[2024] =  12'b000001010111; // 87
storage[2025] =  12'b000000101110; // 46
storage[2026] = -12'b000010110111; // -183
storage[2027] =  12'b000010010000; // 144
storage[2028] =  12'b000011110010; // 242
storage[2029] = -12'b000011110011; // -243
storage[2030] =  12'b000010010011; // 147
storage[2031] =  12'b000001101100; // 108
storage[2032] = -12'b000011110111; // -247
storage[2033] = -12'b000000110100; // -52
storage[2034] =  12'b000010001000; // 136
storage[2035] = -12'b000001011100; // -92
storage[2036] = -12'b000011000010; // -194
storage[2037] =  12'b000010000101; // 133
storage[2038] = -12'b000010010101; // -149
storage[2039] =  12'b000001001101; // 77
storage[2040] =  12'b000011001101; // 205
storage[2041] = -12'b000011101110; // -238
storage[2042] = -12'b000010111101; // -189
storage[2043] = -12'b000000101101; // -45
storage[2044] =  12'b000100110010; // 306
storage[2045] = -12'b000010010110; // -150
storage[2046] = -12'b000001000111; // -71
storage[2047] =  12'b000001101011; // 107
storage[2048] = -12'b000001110011; // -115
storage[2049] = -12'b000001011001; // -89
storage[2050] = -12'b000000110010; // -50
storage[2051] =  12'b000000011010; // 26
storage[2052] = -12'b000011010011; // -211
storage[2053] = -12'b000100111011; // -315
storage[2054] = -12'b000011010010; // -210
storage[2055] = -12'b000001100000; // -96
storage[2056] = -12'b000100110001; // -305
storage[2057] =  12'b000000011010; // 26
storage[2058] =  12'b000010001001; // 137
storage[2059] =  12'b000011000110; // 198
storage[2060] = -12'b000001110011; // -115
storage[2061] = -12'b000001011111; // -95
storage[2062] =  12'b000010011010; // 154
storage[2063] =  12'b000001011010; // 90
storage[2064] = -12'b000101101011; // -363
storage[2065] =  12'b000001011110; // 94
storage[2066] =  12'b000011111101; // 253
storage[2067] =  12'b000000000111; // 7
storage[2068] = -12'b000000101011; // -43
storage[2069] = -12'b000010011110; // -158
storage[2070] = -12'b000001010000; // -80
storage[2071] =  12'b000100000100; // 260
storage[2072] = -12'b000001111101; // -125
storage[2073] = -12'b000100010000; // -272
storage[2074] =  12'b000011000100; // 196
storage[2075] =  12'b000001101001; // 105
storage[2076] = -12'b000010000100; // -132
storage[2077] =  12'b000010100000; // 160
storage[2078] = -12'b000000001010; // -10
storage[2079] =  12'b000010100111; // 167
storage[2080] =  12'b000010111010; // 186
storage[2081] =  12'b000100001001; // 265
storage[2082] = -12'b000000100101; // -37
storage[2083] = -12'b000000111100; // -60
storage[2084] =  12'b000001001110; // 78
storage[2085] =  12'b000010000001; // 129
storage[2086] =  12'b000000000011; // 3
storage[2087] =  12'b000010110011; // 179
storage[2088] =  12'b000101100111; // 359
storage[2089] = -12'b000000110001; // -49
storage[2090] =  12'b000101111010; // 378
storage[2091] =  12'b000100110110; // 310
storage[2092] = -12'b000000010001; // -17
storage[2093] =  12'b000001100100; // 100
storage[2094] =  12'b000111000000; // 448
storage[2095] = -12'b000011110011; // -243
storage[2096] =  12'b000001010111; // 87
storage[2097] =  12'b000010000000; // 128
storage[2098] = -12'b000100001010; // -266
storage[2099] =  12'b000000111010; // 58
storage[2100] =  12'b000000110100; // 52
storage[2101] =  12'b000000011000; // 24
storage[2102] =  12'b000011100101; // 229
storage[2103] =  12'b000000011000; // 24
storage[2104] = -12'b000011010101; // -213
storage[2105] = -12'b000011101000; // -232
storage[2106] = -12'b000001001110; // -78
storage[2107] = -12'b000010111000; // -184
storage[2108] =  12'b000000010110; // 22
storage[2109] =  12'b000000010011; // 19
storage[2110] = -12'b000010101011; // -171
storage[2111] = -12'b000000100110; // -38
storage[2112] =  12'b000000011010; // 26
storage[2113] = -12'b000100010110; // -278
storage[2114] = -12'b001001010001; // -593
storage[2115] =  12'b000000110000; // 48
storage[2116] =  12'b000100001111; // 271
storage[2117] =  12'b000001011010; // 90
storage[2118] =  12'b000011100001; // 225
storage[2119] =  12'b000011110110; // 246
storage[2120] =  12'b000001101011; // 107
storage[2121] =  12'b000011001101; // 205
storage[2122] =  12'b000010100010; // 162
storage[2123] =  12'b000001001011; // 75
storage[2124] = -12'b000001000001; // -65
storage[2125] = -12'b000010010110; // -150
storage[2126] =  12'b000000110001; // 49
storage[2127] =  12'b000001111101; // 125
storage[2128] =  12'b000000111001; // 57
storage[2129] = -12'b000000000010; // -2
storage[2130] = -12'b000001011111; // -95
storage[2131] =  12'b000000100000; // 32
storage[2132] = -12'b000101011010; // -346
storage[2133] =  12'b000001010100; // 84
storage[2134] =  12'b000000101110; // 46
storage[2135] = -12'b000001101100; // -108
storage[2136] = -12'b000000110100; // -52
storage[2137] = -12'b000010010110; // -150
storage[2138] = -12'b000100010100; // -276
storage[2139] =  12'b000001101011; // 107
storage[2140] =  12'b000010011110; // 158
storage[2141] = -12'b000100100101; // -293
storage[2142] = -12'b000011001101; // -205
storage[2143] =  12'b000001010010; // 82
storage[2144] =  12'b000001111001; // 121
storage[2145] = -12'b000000100010; // -34
storage[2146] =  12'b000010100010; // 162
storage[2147] = -12'b000001010100; // -84
storage[2148] = -12'b000100000001; // -257
storage[2149] = -12'b000000011011; // -27
storage[2150] = -12'b000010101101; // -173
storage[2151] = -12'b000101101001; // -361
storage[2152] =  12'b000001100110; // 102
storage[2153] = -12'b000000111011; // -59
storage[2154] =  12'b000100001001; // 265
storage[2155] = -12'b000100001000; // -264
storage[2156] =  12'b000000010011; // 19
storage[2157] =  12'b000000101111; // 47
storage[2158] = -12'b000000100101; // -37
storage[2159] = -12'b000101101100; // -364
storage[2160] = -12'b000100100011; // -291
storage[2161] =  12'b000001001111; // 79
storage[2162] = -12'b000000110101; // -53
storage[2163] = -12'b000011100000; // -224
storage[2164] = -12'b000010101000; // -168
storage[2165] = -12'b000001010110; // -86
storage[2166] = -12'b000000010001; // -17
storage[2167] = -12'b000011000101; // -197
storage[2168] = -12'b000000101011; // -43
storage[2169] =  12'b000110001110; // 398
storage[2170] =  12'b000001001101; // 77
storage[2171] =  12'b000100000101; // 261
storage[2172] = -12'b000001000100; // -68
storage[2173] =  12'b000010111110; // 190
storage[2174] = -12'b000000010001; // -17
storage[2175] = -12'b000000100111; // -39
storage[2176] = -12'b000001010111; // -87
storage[2177] = -12'b000000101111; // -47
storage[2178] =  12'b000000101110; // 46
storage[2179] =  12'b000010000000; // 128
storage[2180] =  12'b000010100110; // 166
storage[2181] = -12'b000000011100; // -28
storage[2182] =  12'b000000011000; // 24
storage[2183] = -12'b000000100011; // -35
storage[2184] = -12'b000000001000; // -8
storage[2185] =  12'b000100101010; // 298
storage[2186] =  12'b000011100100; // 228
storage[2187] =  12'b000111000100; // 452
storage[2188] = -12'b000001000101; // -69
storage[2189] =  12'b000000101101; // 45
storage[2190] = -12'b000010011100; // -156
storage[2191] =  12'b000000000011; // 3
storage[2192] = -12'b000000100001; // -33
storage[2193] =  12'b000010011101; // 157
storage[2194] = -12'b000010101110; // -174
storage[2195] =  12'b000000101000; // 40
storage[2196] = -12'b000000001110; // -14
storage[2197] =  12'b000000100000; // 32
storage[2198] = -12'b000000100000; // -32
storage[2199] =  12'b000010111001; // 185
storage[2200] =  12'b000010100010; // 162
storage[2201] =  12'b000100100001; // 289
storage[2202] =  12'b000011010110; // 214
storage[2203] = -12'b000000010110; // -22
storage[2204] = -12'b000000000110; // -6
storage[2205] =  12'b000010100010; // 162
storage[2206] = -12'b000011111011; // -251
storage[2207] = -12'b000000001000; // -8
storage[2208] = -12'b000010011011; // -155
storage[2209] = -12'b000001101000; // -104
storage[2210] = -12'b000000001001; // -9
storage[2211] =  12'b000000110001; // 49
storage[2212] =  12'b000011011011; // 219
storage[2213] =  12'b000100000101; // 261
storage[2214] =  12'b000101000100; // 324
storage[2215] =  12'b000001000100; // 68
storage[2216] = -12'b000011000000; // -192
storage[2217] = -12'b000011101000; // -232
storage[2218] =  12'b000000110100; // 52
storage[2219] = -12'b000001001000; // -72
storage[2220] = -12'b000011100000; // -224
storage[2221] =  12'b000000010111; // 23
storage[2222] = -12'b000011110101; // -245
storage[2223] =  12'b000001110011; // 115
storage[2224] =  12'b000001110101; // 117
storage[2225] =  12'b000000100111; // 39
storage[2226] =  12'b000000011000; // 24
storage[2227] =  12'b000000100011; // 35
storage[2228] = -12'b000000010000; // -16
storage[2229] =  12'b000000011110; // 30
storage[2230] = -12'b000000110001; // -49
storage[2231] =  12'b000010110001; // 177
storage[2232] =  12'b000001010110; // 86
storage[2233] =  12'b000011000010; // 194
storage[2234] =  12'b000100010111; // 279
storage[2235] =  12'b000010101111; // 175
storage[2236] =  12'b000010100111; // 167
storage[2237] =  12'b000010001110; // 142
storage[2238] =  12'b000100000010; // 258
storage[2239] =  12'b000111011010; // 474
storage[2240] =  12'b000111100111; // 487
storage[2241] =  12'b000000011001; // 25
storage[2242] = -12'b000001011011; // -91
storage[2243] = -12'b000010110101; // -181
storage[2244] = -12'b000000010111; // -23
storage[2245] = -12'b000000001100; // -12
storage[2246] = -12'b000011001111; // -207
storage[2247] =  12'b000001011110; // 94
storage[2248] =  12'b000001111001; // 121
storage[2249] =  12'b000000110010; // 50
storage[2250] = -12'b000000011110; // -30
storage[2251] =  12'b000010110111; // 183
storage[2252] = -12'b000000011110; // -30
storage[2253] = -12'b000011001110; // -206
storage[2254] = -12'b000000011001; // -25
storage[2255] = -12'b000010100100; // -164
storage[2256] = -12'b000100000110; // -262
storage[2257] = -12'b000000111111; // -63
storage[2258] =  12'b000001111010; // 122
storage[2259] =  12'b000100101010; // 298
storage[2260] =  12'b000001000111; // 71
storage[2261] = -12'b000000001000; // -8
storage[2262] =  12'b000001001000; // 72
storage[2263] =  12'b000001110101; // 117
storage[2264] =  12'b000010110010; // 178
storage[2265] =  12'b000100100000; // 288
storage[2266] = -12'b000000001001; // -9
storage[2267] =  12'b000010001010; // 138
storage[2268] = -12'b000000011101; // -29
storage[2269] = -12'b000001111100; // -124
storage[2270] = -12'b000001111110; // -126
storage[2271] =  12'b000001110101; // 117
storage[2272] = -12'b000010000011; // -131
storage[2273] =  12'b000001101000; // 104
storage[2274] =  12'b000010111001; // 185
storage[2275] = -12'b000000010100; // -20
storage[2276] = -12'b000000001001; // -9
storage[2277] =  12'b000000011101; // 29
storage[2278] = -12'b000101010001; // -337
storage[2279] =  12'b000010010000; // 144
storage[2280] =  12'b000000010111; // 23
storage[2281] =  12'b000111001001; // 457
storage[2282] =  12'b000110010000; // 400
storage[2283] = -12'b000000110111; // -55
storage[2284] =  12'b000010011111; // 159
storage[2285] = -12'b000001100001; // -97
storage[2286] = -12'b000000011011; // -27
storage[2287] = -12'b000101011010; // -346
storage[2288] =  12'b000001100001; // 97
storage[2289] =  12'b000001110101; // 117
storage[2290] = -12'b000001011110; // -94
storage[2291] = -12'b000000010110; // -22
storage[2292] =  12'b000001100011; // 99
storage[2293] = -12'b000000011010; // -26
storage[2294] = -12'b000011000101; // -197
storage[2295] = -12'b000001001100; // -76
storage[2296] = -12'b000100011101; // -285
storage[2297] =  12'b000001111011; // 123
storage[2298] = -12'b000100000101; // -261
storage[2299] = -12'b000000011110; // -30
storage[2300] = -12'b000010011010; // -154
storage[2301] = -12'b000001111001; // -121
storage[2302] =  12'b000011001011; // 203
storage[2303] =  12'b000000000100; // 4
storage[2304] =  12'b000011000000; // 192
storage[2305] = -12'b000000101110; // -46
storage[2306] = -12'b000000110010; // -50
storage[2307] = -12'b000011001001; // -201
storage[2308] = -12'b000001100101; // -101
storage[2309] = -12'b000000011001; // -25
storage[2310] =  12'b000000011110; // 30
storage[2311] = -12'b000001010111; // -87
storage[2312] =  12'b000000110110; // 54
storage[2313] = -12'b000011100001; // -225
storage[2314] = -12'b000010110100; // -180
storage[2315] = -12'b000001101111; // -111
storage[2316] =  12'b000011000100; // 196
storage[2317] =  12'b000001101011; // 107
storage[2318] = -12'b000000100001; // -33
storage[2319] = -12'b000000101100; // -44
storage[2320] =  12'b000001110000; // 112
storage[2321] = -12'b000001010010; // -82
storage[2322] = -12'b000000110000; // -48
storage[2323] =  12'b000000110100; // 52
storage[2324] =  12'b000010010101; // 149
storage[2325] =  12'b000011000011; // 195
storage[2326] =  12'b000100000100; // 260
storage[2327] =  12'b000011010011; // 211
storage[2328] = -12'b000001111011; // -123
storage[2329] =  12'b000001101101; // 109
storage[2330] =  12'b000001110100; // 116
storage[2331] =  12'b000010001011; // 139
storage[2332] =  12'b000100001011; // 267
storage[2333] =  12'b000010010001; // 145
storage[2334] =  12'b000001110000; // 112
storage[2335] =  12'b000000000101; // 5
storage[2336] =  12'b000000011110; // 30
storage[2337] = -12'b000000101010; // -42
storage[2338] =  12'b000010001110; // 142
storage[2339] =  12'b000000111010; // 58
storage[2340] = -12'b000000110001; // -49
storage[2341] =  12'b000001010000; // 80
storage[2342] =  12'b000001110111; // 119
storage[2343] =  12'b000010101101; // 173
storage[2344] =  12'b000001010001; // 81
storage[2345] =  12'b000011110100; // 244
storage[2346] = -12'b000000001111; // -15
storage[2347] =  12'b000000101101; // 45
storage[2348] =  12'b000011110110; // 246
storage[2349] =  12'b000010101100; // 172
storage[2350] = -12'b000110100000; // -416
storage[2351] =  12'b000000111100; // 60
storage[2352] =  12'b000001000100; // 68
storage[2353] = -12'b000010100001; // -161
storage[2354] = -12'b000010111001; // -185
storage[2355] =  12'b000001011000; // 88
storage[2356] =  12'b000010110101; // 181
storage[2357] =  12'b000100111000; // 312
storage[2358] = -12'b000000110110; // -54
storage[2359] =  12'b000011100000; // 224
storage[2360] =  12'b000001111001; // 121
storage[2361] = -12'b000000010100; // -20
storage[2362] =  12'b000010110101; // 181
storage[2363] =  12'b000010100011; // 163
storage[2364] = -12'b000000111101; // -61
storage[2365] = -12'b000001111001; // -121
storage[2366] =  12'b000000001101; // 13
storage[2367] = -12'b000010110100; // -180
storage[2368] = -12'b000010100100; // -164
storage[2369] = -12'b000001100110; // -102
storage[2370] =  12'b000000101000; // 40
storage[2371] =  12'b000001111001; // 121
storage[2372] = -12'b000000001010; // -10
storage[2373] =  12'b000001101011; // 107
storage[2374] =  12'b000010100100; // 164
storage[2375] = -12'b000000101111; // -47
storage[2376] = -12'b000000111101; // -61
storage[2377] = -12'b000000111011; // -59
storage[2378] = -12'b000000101011; // -43
storage[2379] =  12'b000011110011; // 243
storage[2380] = -12'b000011101110; // -238
storage[2381] = -12'b000010001011; // -139
storage[2382] =  12'b000011111110; // 254
storage[2383] =  12'b000011110010; // 242
storage[2384] = -12'b000010001100; // -140
storage[2385] =  12'b000101010001; // 337
storage[2386] =  12'b000001100011; // 99
storage[2387] =  12'b000011100101; // 229
storage[2388] = -12'b000000010101; // -21
storage[2389] =  12'b000001010001; // 81
storage[2390] = -12'b000010110001; // -177
storage[2391] = -12'b000011111001; // -249
storage[2392] =  12'b000001100001; // 97
storage[2393] =  12'b000000011100; // 28
storage[2394] = -12'b000000111101; // -61
storage[2395] = -12'b000100110000; // -304
storage[2396] = -12'b000010110010; // -178
storage[2397] =  12'b000010000000; // 128
storage[2398] = -12'b000111011101; // -477
storage[2399] = -12'b000101100011; // -355
storage[2400] = -12'b000010111111; // -191
storage[2401] =  12'b000001001101; // 77
storage[2402] = -12'b000001011111; // -95
storage[2403] = -12'b000000000010; // -2
storage[2404] =  12'b000000101101; // 45
storage[2405] = -12'b000001101110; // -110
storage[2406] = -12'b000010001010; // -138
storage[2407] = -12'b000000011010; // -26
storage[2408] = -12'b000011001001; // -201
storage[2409] = -12'b000011101100; // -236
storage[2410] = -12'b000011000110; // -198
storage[2411] = -12'b000010011101; // -157
storage[2412] = -12'b000011101011; // -235
storage[2413] = -12'b000001000100; // -68
storage[2414] = -12'b000000010001; // -17
storage[2415] =  12'b000100011010; // 282
storage[2416] =  12'b000000010000; // 16
storage[2417] =  12'b000000001011; // 11
storage[2418] =  12'b000001010000; // 80
storage[2419] =  12'b000001010110; // 86
storage[2420] =  12'b000011110110; // 246
storage[2421] =  12'b000011100100; // 228
storage[2422] =  12'b000001100001; // 97
storage[2423] =  12'b000110011010; // 410
storage[2424] =  12'b000010101111; // 175
storage[2425] =  12'b000001011101; // 93
storage[2426] =  12'b000100101011; // 299
storage[2427] =  12'b000010101101; // 173
storage[2428] =  12'b000010010111; // 151
storage[2429] =  12'b000010110111; // 183
storage[2430] =  12'b000100100011; // 291
storage[2431] =  12'b000011000100; // 196
storage[2432] =  12'b000010100100; // 164
storage[2433] =  12'b000100001000; // 264
storage[2434] = -12'b000001001100; // -76
storage[2435] =  12'b000001100001; // 97
storage[2436] =  12'b000010001110; // 142
storage[2437] =  12'b000000101100; // 44
storage[2438] = -12'b000000101100; // -44
storage[2439] =  12'b000100001111; // 271
storage[2440] =  12'b000110111101; // 445
storage[2441] =  12'b000010111100; // 188
storage[2442] =  12'b000100100101; // 293
storage[2443] =  12'b000100100000; // 288
storage[2444] =  12'b000001101111; // 111
storage[2445] = -12'b000001010101; // -85
storage[2446] =  12'b000001101010; // 106
storage[2447] =  12'b000000011010; // 26
storage[2448] =  12'b000010000110; // 134
storage[2449] = -12'b000000011011; // -27
storage[2450] = -12'b000011001000; // -200
storage[2451] = -12'b000011101100; // -236
storage[2452] =  12'b000010101100; // 172
storage[2453] = -12'b000000101101; // -45
storage[2454] = -12'b000010000101; // -133
storage[2455] =  12'b000110111111; // 447
storage[2456] =  12'b000001111011; // 123
storage[2457] = -12'b000001111010; // -122
storage[2458] =  12'b000000110001; // 49
storage[2459] =  12'b000000010110; // 22
storage[2460] =  12'b000100011001; // 281
storage[2461] = -12'b000100011010; // -282
storage[2462] = -12'b000000111010; // -58
storage[2463] =  12'b000000001011; // 11
storage[2464] = -12'b000000001000; // -8
storage[2465] =  12'b000011011100; // 220
storage[2466] = -12'b000010010011; // -147
storage[2467] = -12'b000011010110; // -214
storage[2468] =  12'b000000100111; // 39
storage[2469] =  12'b000010001011; // 139
storage[2470] = -12'b000010011001; // -153
storage[2471] = -12'b000000011110; // -30
storage[2472] = -12'b000010011000; // -152
storage[2473] =  12'b000000100100; // 36
storage[2474] = -12'b000011101000; // -232
storage[2475] = -12'b000011010010; // -210
storage[2476] = -12'b000000111000; // -56
storage[2477] =  12'b000010000000; // 128
storage[2478] = -12'b000011110001; // -241
storage[2479] = -12'b000000000001; // -1
storage[2480] =  12'b000001001011; // 75
storage[2481] = -12'b000001000010; // -66
storage[2482] = -12'b001000001010; // -522
storage[2483] = -12'b000010010111; // -151
storage[2484] = -12'b000001001101; // -77
storage[2485] = -12'b000000101010; // -42
storage[2486] =  12'b000000001100; // 12
storage[2487] = -12'b000010000111; // -135
storage[2488] =  12'b000000111110; // 62
storage[2489] =  12'b000101111101; // 381
storage[2490] =  12'b000001011010; // 90
storage[2491] = -12'b000100010000; // -272
storage[2492] =  12'b000000111000; // 56
storage[2493] = -12'b000000000010; // -2
storage[2494] =  12'b000010000100; // 132
storage[2495] =  12'b000011111001; // 249
storage[2496] = -12'b000010000101; // -133
storage[2497] = -12'b000001111000; // -120
storage[2498] =  12'b000000001000; // 8
storage[2499] =  12'b000001010100; // 84
storage[2500] =  12'b000010101000; // 168
storage[2501] =  12'b000001000001; // 65
storage[2502] = -12'b000000001101; // -13
storage[2503] =  12'b000010000001; // 129
storage[2504] =  12'b000000101101; // 45
storage[2505] = -12'b000001110100; // -116
storage[2506] = -12'b000000110110; // -54
storage[2507] = -12'b000000100111; // -39
storage[2508] =  12'b000100101110; // 302
storage[2509] = -12'b001000110110; // -566
storage[2510] = -12'b000010010000; // -144
storage[2511] =  12'b000011111010; // 250
storage[2512] =  12'b000001111101; // 125
storage[2513] =  12'b000001001110; // 78
storage[2514] =  12'b000001001001; // 73
storage[2515] = -12'b000010110110; // -182
storage[2516] = -12'b000010111011; // -187
storage[2517] = -12'b000001001111; // -79
storage[2518] = -12'b000110101100; // -428
storage[2519] = -12'b000001001111; // -79
storage[2520] = -12'b000011000100; // -196
storage[2521] =  12'b000011010001; // 209
storage[2522] =  12'b000010000110; // 134
storage[2523] =  12'b000010010011; // 147
storage[2524] =  12'b000000111001; // 57
storage[2525] =  12'b000011000011; // 195
storage[2526] = -12'b000010011111; // -159
storage[2527] =  12'b000000000110; // 6
storage[2528] = -12'b000110010010; // -402
storage[2529] = -12'b001001010110; // -598
storage[2530] = -12'b000001000010; // -66
storage[2531] = -12'b000001110100; // -116
storage[2532] =  12'b000011000010; // 194
storage[2533] =  12'b000010110101; // 181
storage[2534] = -12'b000001010101; // -85
storage[2535] = -12'b000100000110; // -262
storage[2536] =  12'b000011100001; // 225
storage[2537] =  12'b000010101100; // 172
storage[2538] = -12'b000010100000; // -160
storage[2539] =  12'b000001001000; // 72
storage[2540] =  12'b000010101010; // 170
storage[2541] =  12'b000100101011; // 299
storage[2542] =  12'b000100100000; // 288
storage[2543] = -12'b000010100010; // -162
storage[2544] = -12'b000001100011; // -99
storage[2545] =  12'b000101001011; // 331
storage[2546] =  12'b000100011011; // 283
storage[2547] = -12'b000001100100; // -100
storage[2548] =  12'b000010111010; // 186
storage[2549] =  12'b000101001110; // 334
storage[2550] =  12'b000000000111; // 7
storage[2551] = -12'b000000011010; // -26
storage[2552] = -12'b000000000010; // -2
storage[2553] = -12'b000100001010; // -266
storage[2554] = -12'b000000111111; // -63
storage[2555] = -12'b000011101001; // -233
storage[2556] = -12'b000101001000; // -328
storage[2557] =  12'b000001111010; // 122
storage[2558] =  12'b000001110101; // 117
storage[2559] =  12'b000101000001; // 321
storage[2560] = -12'b000001000010; // -66
storage[2561] = -12'b000011010110; // -214
storage[2562] = -12'b000100100110; // -294
storage[2563] = -12'b001010100101; // -677
storage[2564] = -12'b001000100000; // -544
storage[2565] = -12'b000001011000; // -88
storage[2566] =  12'b000001011011; // 91
storage[2567] =  12'b000111101010; // 490
storage[2568] =  12'b000010001000; // 136
storage[2569] =  12'b000100100001; // 289
storage[2570] =  12'b000101101001; // 361
storage[2571] =  12'b000000111010; // 58
storage[2572] =  12'b000100011101; // 285
storage[2573] =  12'b000110010101; // 405
storage[2574] =  12'b000011000110; // 198
storage[2575] =  12'b000011000001; // 193
storage[2576] = -12'b000001000000; // -64
storage[2577] =  12'b000011110001; // 241
storage[2578] = -12'b000000001010; // -10
storage[2579] =  12'b000001110110; // 118
storage[2580] =  12'b000000110010; // 50
storage[2581] =  12'b000001000100; // 68
storage[2582] = -12'b000001000110; // -70
storage[2583] =  12'b000010011011; // 155
storage[2584] =  12'b000010000100; // 132
storage[2585] =  12'b000100000101; // 261
storage[2586] = -12'b000001101001; // -105
storage[2587] =  12'b000000111100; // 60
storage[2588] = -12'b000001101011; // -107
storage[2589] = -12'b000010010110; // -150
storage[2590] = -12'b000000001101; // -13
storage[2591] = -12'b000001100001; // -97
storage[2592] = -12'b000010111001; // -185
storage[2593] =  12'b000000100000; // 32
storage[2594] =  12'b000000010000; // 16
storage[2595] = -12'b000010101001; // -169
storage[2596] = -12'b000010011110; // -158
storage[2597] = -12'b000001100011; // -99
storage[2598] = -12'b000110101100; // -428
storage[2599] =  12'b000001011100; // 92
storage[2600] =  12'b000010000000; // 128
storage[2601] = -12'b000110110011; // -435
storage[2602] = -12'b000101000111; // -327
storage[2603] = -12'b000000111000; // -56
storage[2604] =  12'b000001000000; // 64
storage[2605] = -12'b000010101110; // -174
storage[2606] = -12'b000010110001; // -177
storage[2607] =  12'b000010011001; // 153
storage[2608] = -12'b000000110011; // -51
storage[2609] = -12'b000001101100; // -108
storage[2610] =  12'b000000010001; // 17
storage[2611] = -12'b000001100110; // -102
storage[2612] =  12'b000000101001; // 41
storage[2613] =  12'b000011001100; // 204
storage[2614] =  12'b000000110001; // 49
storage[2615] =  12'b000110101110; // 430
storage[2616] =  12'b000101000110; // 326
storage[2617] =  12'b000100101010; // 298
storage[2618] =  12'b000110001110; // 398
storage[2619] =  12'b000011111100; // 252
storage[2620] = -12'b000010100111; // -167
storage[2621] = -12'b000101000000; // -320
storage[2622] = -12'b000001110110; // -118
storage[2623] = -12'b000001110011; // -115
storage[2624] = -12'b000001011101; // -93
storage[2625] =  12'b000010111110; // 190
storage[2626] =  12'b000010011110; // 158
storage[2627] =  12'b000001010001; // 81
storage[2628] =  12'b000010111011; // 187
storage[2629] =  12'b000010000011; // 131
storage[2630] =  12'b000001110000; // 112
storage[2631] = -12'b000010100111; // -167
storage[2632] = -12'b000001110110; // -118
storage[2633] = -12'b000000000111; // -7
storage[2634] =  12'b000001010010; // 82
storage[2635] = -12'b000011000100; // -196
storage[2636] =  12'b000000110000; // 48
storage[2637] =  12'b000011011011; // 219
storage[2638] = -12'b000000111000; // -56
storage[2639] = -12'b000101110010; // -370
storage[2640] = -12'b000000100000; // -32
storage[2641] =  12'b000111010010; // 466
storage[2642] =  12'b000010101101; // 173
storage[2643] = -12'b000100000000; // -256
storage[2644] =  12'b000100001000; // 264
storage[2645] =  12'b000100011100; // 284
storage[2646] =  12'b000000100010; // 34
storage[2647] = -12'b000010010111; // -151
storage[2648] = -12'b000011101010; // -234
storage[2649] = -12'b000010010001; // -145
storage[2650] =  12'b000101011010; // 346
storage[2651] =  12'b000101000111; // 327
storage[2652] = -12'b000010110100; // -180
storage[2653] =  12'b000010101111; // 175
storage[2654] =  12'b000011000110; // 198
storage[2655] =  12'b000010010001; // 145
storage[2656] =  12'b000010010110; // 150
storage[2657] =  12'b000010110011; // 179
storage[2658] = -12'b000000000001; // -1
storage[2659] =  12'b000101101111; // 367
storage[2660] =  12'b000011101001; // 233
storage[2661] = -12'b000000001001; // -9
storage[2662] = -12'b000100001101; // -269
storage[2663] = -12'b000010110001; // -177
storage[2664] = -12'b000001000101; // -69
storage[2665] =  12'b000010110000; // 176
storage[2666] = -12'b000000110100; // -52
storage[2667] =  12'b000010101000; // 168
storage[2668] = -12'b000100100010; // -290
storage[2669] =  12'b000001101011; // 107
storage[2670] =  12'b000011001101; // 205
storage[2671] = -12'b000000010111; // -23
storage[2672] =  12'b000010000011; // 131
storage[2673] = -12'b000000110001; // -49
storage[2674] =  12'b000000110110; // 54
storage[2675] = -12'b000001001001; // -73
storage[2676] =  12'b000010110110; // 182
storage[2677] = -12'b000001111111; // -127
storage[2678] = -12'b000000010100; // -20
storage[2679] = -12'b000011010010; // -210
storage[2680] = -12'b000001011101; // -93
storage[2681] =  12'b000011001111; // 207
storage[2682] =  12'b000110101001; // 425
storage[2683] = -12'b000011111011; // -251
storage[2684] = -12'b000011010011; // -211
storage[2685] = -12'b000001011000; // -88
storage[2686] =  12'b000000101111; // 47
storage[2687] =  12'b000010010010; // 146
storage[2688] = -12'b000101001111; // -335
storage[2689] = -12'b000000010111; // -23
storage[2690] =  12'b000001011011; // 91
storage[2691] = -12'b000010011011; // -155
storage[2692] = -12'b000101100001; // -353
storage[2693] =  12'b000001110110; // 118
storage[2694] =  12'b000001101111; // 111
storage[2695] = -12'b000001000000; // -64
storage[2696] = -12'b000000110010; // -50
storage[2697] =  12'b000001010001; // 81
storage[2698] =  12'b000010111001; // 185
storage[2699] = -12'b000000011101; // -29
storage[2700] = -12'b000100110010; // -306
storage[2701] =  12'b000000101111; // 47
storage[2702] =  12'b000011011001; // 217
storage[2703] =  12'b000100101010; // 298
storage[2704] =  12'b000010010010; // 146
storage[2705] =  12'b000100111110; // 318
storage[2706] =  12'b000000100101; // 37
storage[2707] =  12'b000010100110; // 166
storage[2708] = -12'b000010000101; // -133
storage[2709] = -12'b000001011111; // -95
storage[2710] = -12'b000001001001; // -73
storage[2711] = -12'b000001111110; // -126
storage[2712] = -12'b000010110011; // -179
storage[2713] =  12'b000010010011; // 147
storage[2714] =  12'b000011010010; // 210
storage[2715] =  12'b000101111000; // 376
storage[2716] =  12'b000001011101; // 93
storage[2717] =  12'b000000101100; // 44
storage[2718] =  12'b000101110101; // 373
storage[2719] =  12'b000010000110; // 134
storage[2720] = -12'b000000101010; // -42
storage[2721] = -12'b000011011011; // -219
storage[2722] =  12'b000000111111; // 63
storage[2723] = -12'b000010101001; // -169
storage[2724] =  12'b000011011010; // 218
storage[2725] =  12'b000000010010; // 18
storage[2726] = -12'b000001001000; // -72
storage[2727] = -12'b000101011111; // -351
storage[2728] = -12'b000000110001; // -49
storage[2729] = -12'b000001111010; // -122
storage[2730] = -12'b000100100010; // -290
storage[2731] = -12'b000010010110; // -150
storage[2732] =  12'b000001010011; // 83
storage[2733] =  12'b000011111100; // 252
storage[2734] =  12'b000100000010; // 258
storage[2735] =  12'b000011001111; // 207
storage[2736] =  12'b000001101110; // 110
storage[2737] = -12'b000001000010; // -66
storage[2738] =  12'b000010011001; // 153
storage[2739] =  12'b000001000111; // 71
storage[2740] = -12'b000001101100; // -108
storage[2741] =  12'b000010111001; // 185
storage[2742] = -12'b000010000010; // -130
storage[2743] = -12'b000010001001; // -137
storage[2744] =  12'b000010001101; // 141
storage[2745] =  12'b000010101000; // 168
storage[2746] = -12'b000000110100; // -52
storage[2747] =  12'b000001100110; // 102
storage[2748] =  12'b000111010000; // 464
storage[2749] =  12'b000010000101; // 133
storage[2750] = -12'b000000111011; // -59
storage[2751] = -12'b000010000011; // -131
storage[2752] = -12'b000010111000; // -184
storage[2753] = -12'b000000010110; // -22
storage[2754] =  12'b000010100011; // 163
storage[2755] =  12'b000001110000; // 112
storage[2756] = -12'b000001100100; // -100
storage[2757] = -12'b000001000001; // -65
storage[2758] = -12'b000000110100; // -52
storage[2759] = -12'b000011010100; // -212
storage[2760] = -12'b000010000111; // -135
storage[2761] = -12'b000011010000; // -208
storage[2762] = -12'b000010011000; // -152
storage[2763] =  12'b000011100010; // 226
storage[2764] =  12'b000011001111; // 207
storage[2765] =  12'b000100111000; // 312
storage[2766] = -12'b000000100100; // -36
storage[2767] =  12'b000011100001; // 225
storage[2768] = -12'b000000101100; // -44
storage[2769] = -12'b000010101100; // -172
storage[2770] =  12'b000000011101; // 29
storage[2771] =  12'b000100100010; // 290
storage[2772] =  12'b000001111000; // 120
storage[2773] =  12'b000011000101; // 197
storage[2774] = -12'b000010000010; // -130
storage[2775] = -12'b000010100001; // -161
storage[2776] =  12'b000010110000; // 176
storage[2777] = -12'b000101110111; // -375
storage[2778] = -12'b000111011100; // -476
storage[2779] = -12'b000010000010; // -130
storage[2780] = -12'b000011110101; // -245
storage[2781] = -12'b000001111010; // -122
storage[2782] = -12'b000110010000; // -400
storage[2783] = -12'b000011010110; // -214
storage[2784] =  12'b000010011010; // 154
storage[2785] = -12'b000010111100; // -188
storage[2786] =  12'b000000100011; // 35
storage[2787] =  12'b000001000001; // 65
storage[2788] =  12'b000000111011; // 59
storage[2789] = -12'b000000101011; // -43
storage[2790] = -12'b000011011000; // -216
storage[2791] = -12'b000100010111; // -279
storage[2792] = -12'b000000001000; // -8
storage[2793] = -12'b000001011111; // -95
storage[2794] = -12'b000001010101; // -85
storage[2795] =  12'b000011110001; // 241
storage[2796] = -12'b000010110000; // -176
storage[2797] =  12'b000010110010; // 178
storage[2798] =  12'b000110101001; // 425
storage[2799] = -12'b000000010011; // -19
storage[2800] = -12'b000000000110; // -6
storage[2801] =  12'b000000101001; // 41
storage[2802] =  12'b000000001100; // 12
storage[2803] =  12'b000010000110; // 134
storage[2804] =  12'b000000111100; // 60
storage[2805] =  12'b000001101010; // 106
storage[2806] =  12'b000000000110; // 6
storage[2807] = -12'b000001111011; // -123
storage[2808] =  12'b000000101000; // 40
storage[2809] =  12'b000010100001; // 161
storage[2810] =  12'b000000000001; // 1
storage[2811] = -12'b000101011000; // -344
storage[2812] =  12'b000001011001; // 89
storage[2813] = -12'b000010000101; // -133
storage[2814] = -12'b000000010010; // -18
storage[2815] = -12'b000011101010; // -234
storage[2816] = -12'b000101100001; // -353
storage[2817] = -12'b000001000111; // -71
storage[2818] = -12'b000001011111; // -95
storage[2819] = -12'b000001100111; // -103
storage[2820] = -12'b000010010001; // -145
storage[2821] = -12'b000001010000; // -80
storage[2822] =  12'b000000111011; // 59
storage[2823] =  12'b000000010111; // 23
storage[2824] =  12'b000011011011; // 219
storage[2825] =  12'b000101001001; // 329
storage[2826] =  12'b000101110010; // 370
storage[2827] = -12'b000000100110; // -38
storage[2828] =  12'b000000011010; // 26
storage[2829] = -12'b000000010011; // -19
storage[2830] =  12'b000010100011; // 163
storage[2831] =  12'b000011101110; // 238
storage[2832] =  12'b000101000101; // 325
storage[2833] =  12'b000001101010; // 106
storage[2834] =  12'b000010101111; // 175
storage[2835] =  12'b000010010101; // 149
storage[2836] =  12'b000000100010; // 34
storage[2837] =  12'b000000110011; // 51
storage[2838] =  12'b000101101111; // 367
storage[2839] = -12'b000000101011; // -43
storage[2840] =  12'b000011010100; // 212
storage[2841] =  12'b000101001100; // 332
storage[2842] =  12'b000000101011; // 43
storage[2843] = -12'b000001101110; // -110
storage[2844] = -12'b000001100110; // -102
storage[2845] = -12'b000000000110; // -6
storage[2846] = -12'b000000110010; // -50
storage[2847] = -12'b000000011001; // -25
storage[2848] =  12'b000010000010; // 130
storage[2849] =  12'b000010110011; // 179
storage[2850] = -12'b000100001111; // -271
storage[2851] =  12'b000001000000; // 64
storage[2852] =  12'b000000101100; // 44
storage[2853] = -12'b000101100001; // -353
storage[2854] = -12'b000100001000; // -264
storage[2855] = -12'b000001001001; // -73
storage[2856] = -12'b000001011111; // -95
storage[2857] = -12'b000011100010; // -226
storage[2858] =  12'b000001101011; // 107
storage[2859] = -12'b000001111110; // -126
storage[2860] = -12'b000110110010; // -434
storage[2861] = -12'b001000001000; // -520
storage[2862] = -12'b001001011110; // -606
storage[2863] = -12'b000001011111; // -95
storage[2864] =  12'b000011010100; // 212
storage[2865] =  12'b000000110101; // 53
storage[2866] = -12'b000000100110; // -38
storage[2867] =  12'b000010110111; // 183
storage[2868] =  12'b000000110100; // 52
storage[2869] = -12'b000101101010; // -362
storage[2870] = -12'b000001111100; // -124
storage[2871] = -12'b000111010000; // -464
storage[2872] = -12'b000010011100; // -156
storage[2873] =  12'b000000001011; // 11
storage[2874] =  12'b000001001101; // 77
storage[2875] = -12'b000000111100; // -60
storage[2876] =  12'b000011110111; // 247
storage[2877] =  12'b000011101000; // 232
storage[2878] = -12'b000011000001; // -193
storage[2879] = -12'b000110101001; // -425
storage[2880] = -12'b000101110000; // -368
storage[2881] =  12'b000010010100; // 148
storage[2882] = -12'b000000110011; // -51
storage[2883] = -12'b000011001000; // -200
storage[2884] =  12'b000010000011; // 131
storage[2885] =  12'b000100000010; // 258
storage[2886] = -12'b000001100110; // -102
storage[2887] =  12'b000100110000; // 304
storage[2888] =  12'b000001011110; // 94
storage[2889] =  12'b000010010000; // 144
storage[2890] =  12'b000000000010; // 2
storage[2891] =  12'b000000011011; // 27
storage[2892] =  12'b000011010010; // 210
storage[2893] = -12'b000000001011; // -11
storage[2894] = -12'b000001000101; // -69
storage[2895] =  12'b000000110110; // 54
storage[2896] =  12'b000001110100; // 116
storage[2897] = -12'b000010010000; // -144
storage[2898] =  12'b000000101101; // 45
storage[2899] = -12'b000001111101; // -125
storage[2900] =  12'b000100000111; // 263
storage[2901] =  12'b000011000101; // 197
storage[2902] =  12'b000010100101; // 165
storage[2903] =  12'b000000011101; // 29
storage[2904] =  12'b000000111100; // 60
storage[2905] = -12'b000000110110; // -54
storage[2906] = -12'b000000010001; // -17
storage[2907] =  12'b000100000111; // 263
storage[2908] = -12'b000011110011; // -243
storage[2909] = -12'b000000101011; // -43
storage[2910] = -12'b000010001011; // -139
storage[2911] = -12'b000000110010; // -50
storage[2912] = -12'b000100101001; // -297
storage[2913] =  12'b000011000000; // 192
storage[2914] = -12'b000001111000; // -120
storage[2915] = -12'b000000010010; // -18
storage[2916] =  12'b000010111010; // 186
storage[2917] = -12'b000001001110; // -78
storage[2918] = -12'b000000011110; // -30
storage[2919] =  12'b000010101101; // 173
storage[2920] =  12'b000001001010; // 74
storage[2921] =  12'b000001111111; // 127
storage[2922] =  12'b000001100000; // 96
storage[2923] =  12'b000001100100; // 100
storage[2924] = -12'b000001111011; // -123
storage[2925] =  12'b000001111011; // 123
storage[2926] =  12'b000001011110; // 94
storage[2927] =  12'b000011000001; // 193
storage[2928] = -12'b000010010011; // -147
storage[2929] =  12'b000100011010; // 282
storage[2930] =  12'b000010000010; // 130
storage[2931] = -12'b000010111111; // -191
storage[2932] =  12'b000111011111; // 479
storage[2933] = -12'b000000110111; // -55
storage[2934] =  12'b000000011000; // 24
storage[2935] = -12'b000000011011; // -27
storage[2936] =  12'b000010000010; // 130
storage[2937] =  12'b000000011000; // 24
storage[2938] = -12'b000000001110; // -14
storage[2939] =  12'b000000000100; // 4
storage[2940] =  12'b000010101100; // 172
storage[2941] =  12'b000000010111; // 23
storage[2942] =  12'b000010001101; // 141
storage[2943] =  12'b000000001101; // 13
storage[2944] = -12'b000001110111; // -119
storage[2945] = -12'b000001000110; // -70
storage[2946] =  12'b000100101111; // 303
storage[2947] =  12'b000000101111; // 47
storage[2948] = -12'b000011100000; // -224
storage[2949] =  12'b000001100100; // 100
storage[2950] = -12'b000010001001; // -137
storage[2951] = -12'b000001011001; // -89
storage[2952] =  12'b000001000111; // 71
storage[2953] =  12'b000001101001; // 105
storage[2954] = -12'b000001010111; // -87
storage[2955] =  12'b000001010001; // 81
storage[2956] =  12'b000001110010; // 114
storage[2957] =  12'b000001100001; // 97
storage[2958] = -12'b000010010110; // -150
storage[2959] =  12'b000000111001; // 57
storage[2960] =  12'b000100111100; // 316
storage[2961] =  12'b000001101011; // 107
storage[2962] = -12'b000000001101; // -13
storage[2963] = -12'b000010101110; // -174
storage[2964] = -12'b000110100100; // -420
storage[2965] = -12'b000001111100; // -124
storage[2966] = -12'b000110011000; // -408
storage[2967] = -12'b000100100011; // -291
storage[2968] =  12'b000100111010; // 314
storage[2969] =  12'b000101001001; // 329
storage[2970] =  12'b000110111101; // 445
storage[2971] =  12'b000001001111; // 79
storage[2972] = -12'b000100111000; // -312
storage[2973] = -12'b000011010010; // -210
storage[2974] =  12'b000000100100; // 36
storage[2975] = -12'b000101000001; // -321
storage[2976] = -12'b000110001011; // -395
storage[2977] =  12'b000110101010; // 426
storage[2978] =  12'b000001101100; // 108
storage[2979] = -12'b000000001001; // -9
storage[2980] =  12'b000010101100; // 172
storage[2981] = -12'b000001001101; // -77
storage[2982] =  12'b000010000101; // 133
storage[2983] = -12'b000001001010; // -74
storage[2984] = -12'b000001110110; // -118
storage[2985] =  12'b000001000000; // 64
storage[2986] = -12'b000010001010; // -138
storage[2987] = -12'b000101100011; // -355
storage[2988] = -12'b000010111011; // -187
storage[2989] =  12'b000000110101; // 53
storage[2990] =  12'b000010110010; // 178
storage[2991] = -12'b000010100000; // -160
storage[2992] = -12'b000011000100; // -196
storage[2993] = -12'b000001111101; // -125
storage[2994] =  12'b000001011010; // 90
storage[2995] =  12'b000000010111; // 23
storage[2996] =  12'b000010101001; // 169
storage[2997] =  12'b000000111001; // 57
storage[2998] = -12'b000101001000; // -328
storage[2999] = -12'b000011000011; // -195
storage[3000] = -12'b000000101100; // -44
storage[3001] = -12'b000001011100; // -92
storage[3002] = -12'b000011011100; // -220
storage[3003] = -12'b000011101110; // -238
storage[3004] = -12'b000011000010; // -194
storage[3005] = -12'b000001010001; // -81
storage[3006] = -12'b000001011100; // -92
storage[3007] =  12'b000001011111; // 95
storage[3008] =  12'b000010101110; // 174
storage[3009] =  12'b000001101100; // 108
storage[3010] =  12'b000001011101; // 93
storage[3011] =  12'b000100111110; // 318
storage[3012] =  12'b000001010011; // 83
storage[3013] = -12'b000001100010; // -98
storage[3014] =  12'b000000001001; // 9
storage[3015] = -12'b000000110101; // -53
storage[3016] = -12'b000010000001; // -129
storage[3017] = -12'b000100111111; // -319
storage[3018] = -12'b001000011010; // -538
storage[3019] =  12'b000001101101; // 109
storage[3020] =  12'b000000111010; // 58
storage[3021] = -12'b000010101101; // -173
storage[3022] =  12'b000001000010; // 66
storage[3023] =  12'b000011100100; // 228
storage[3024] = -12'b000000110111; // -55
storage[3025] = -12'b000010100110; // -166
storage[3026] = -12'b000001100000; // -96
storage[3027] = -12'b000011011110; // -222
storage[3028] = -12'b000001001000; // -72
storage[3029] =  12'b000010000110; // 134
storage[3030] =  12'b000001001111; // 79
storage[3031] =  12'b000001111100; // 124
storage[3032] =  12'b000000111011; // 59
storage[3033] =  12'b000000101111; // 47
storage[3034] =  12'b000000100011; // 35
storage[3035] = -12'b000000100011; // -35
storage[3036] =  12'b000011011110; // 222
storage[3037] =  12'b000001011110; // 94
storage[3038] =  12'b000001100110; // 102
storage[3039] =  12'b000001010101; // 85
storage[3040] =  12'b000011111000; // 248
storage[3041] =  12'b000010110111; // 183
storage[3042] =  12'b000010001010; // 138
storage[3043] = -12'b000101111010; // -378
storage[3044] = -12'b000010110010; // -178
storage[3045] = -12'b000000000110; // -6
storage[3046] = -12'b001101101000; // -872
storage[3047] = -12'b000101110011; // -371
storage[3048] = -12'b000100100000; // -288
storage[3049] = -12'b000010101110; // -174
storage[3050] =  12'b000001010000; // 80
storage[3051] = -12'b000010010111; // -151
storage[3052] =  12'b000000010011; // 19
storage[3053] =  12'b000001100010; // 98
storage[3054] = -12'b000001001111; // -79
storage[3055] = -12'b000001111111; // -127
storage[3056] = -12'b000100001100; // -268
storage[3057] = -12'b000010000101; // -133
storage[3058] = -12'b000010110111; // -183
storage[3059] = -12'b000000100100; // -36
storage[3060] =  12'b000001111100; // 124
storage[3061] = -12'b000001011010; // -90
storage[3062] =  12'b000010111001; // 185
storage[3063] =  12'b000011010010; // 210
storage[3064] = -12'b000000000001; // -1
storage[3065] = -12'b000001111111; // -127
storage[3066] =  12'b000000010100; // 20
storage[3067] =  12'b000010110010; // 178
storage[3068] = -12'b000000100011; // -35
storage[3069] =  12'b000011100000; // 224
storage[3070] = -12'b000000111010; // -58
storage[3071] = -12'b000010000000; // -128
storage[3072] = -12'b000010000110; // -134
storage[3073] = -12'b000001110110; // -118
storage[3074] =  12'b000001000101; // 69
storage[3075] =  12'b000011110100; // 244
storage[3076] =  12'b000011000000; // 192
storage[3077] =  12'b000001100111; // 103
storage[3078] =  12'b000101000111; // 327
storage[3079] =  12'b000011000001; // 193
storage[3080] = -12'b000001000101; // -69
storage[3081] = -12'b000000010011; // -19
storage[3082] = -12'b000011000111; // -199
storage[3083] = -12'b000010001100; // -140
storage[3084] = -12'b000000111000; // -56
storage[3085] = -12'b000000110100; // -52
storage[3086] = -12'b000011111111; // -255
storage[3087] =  12'b000001011011; // 91
storage[3088] = -12'b000011001101; // -205
storage[3089] = -12'b000001001011; // -75
storage[3090] = -12'b000010010001; // -145
storage[3091] = -12'b000010111011; // -187
storage[3092] =  12'b000001100101; // 101
storage[3093] =  12'b000001000001; // 65
storage[3094] = -12'b000010010000; // -144
storage[3095] =  12'b000001010011; // 83
storage[3096] =  12'b000001110010; // 114
storage[3097] =  12'b000010001101; // 141
storage[3098] = -12'b000011110000; // -240
storage[3099] = -12'b000111101000; // -488
storage[3100] =  12'b000011011001; // 217
storage[3101] =  12'b000001100000; // 96
storage[3102] =  12'b000000111010; // 58
storage[3103] = -12'b000000100101; // -37
storage[3104] = -12'b000010001111; // -143
storage[3105] = -12'b000000011000; // -24
storage[3106] =  12'b000001010110; // 86
storage[3107] = -12'b000010011111; // -159
storage[3108] =  12'b000001111101; // 125
storage[3109] = -12'b000000100010; // -34
storage[3110] = -12'b000111100110; // -486
storage[3111] = -12'b000100100110; // -294
storage[3112] =  12'b000000110101; // 53
storage[3113] = -12'b000001000010; // -66
storage[3114] = -12'b000011010010; // -210
storage[3115] = -12'b000010100000; // -160
storage[3116] = -12'b000000101001; // -41
storage[3117] = -12'b000000100111; // -39
storage[3118] =  12'b000011101101; // 237
storage[3119] = -12'b000000001011; // -11
storage[3120] =  12'b000001011111; // 95
storage[3121] = -12'b000100011111; // -287
storage[3122] = -12'b000001100111; // -103
storage[3123] =  12'b000001011010; // 90
storage[3124] =  12'b000011010111; // 215
storage[3125] = -12'b000000011000; // -24
storage[3126] =  12'b000001011010; // 90
storage[3127] =  12'b000011111110; // 254
storage[3128] =  12'b000001010011; // 83
storage[3129] =  12'b000000010011; // 19
storage[3130] =  12'b000001010001; // 81
storage[3131] =  12'b000001110110; // 118
storage[3132] =  12'b000011010100; // 212
storage[3133] = -12'b000000001100; // -12
storage[3134] =  12'b000000000001; // 1
storage[3135] =  12'b000001111100; // 124
storage[3136] =  12'b000010001001; // 137
storage[3137] =  12'b000001001101; // 77
storage[3138] = -12'b000011001000; // -200
storage[3139] = -12'b000001101110; // -110
storage[3140] = -12'b000001101010; // -106
storage[3141] = -12'b000001101011; // -107
storage[3142] = -12'b000000100100; // -36
storage[3143] = -12'b000001000101; // -69
storage[3144] = -12'b000011101010; // -234
storage[3145] =  12'b000100100110; // 294
storage[3146] =  12'b000101111101; // 381
storage[3147] =  12'b000000100100; // 36
storage[3148] = -12'b000100000010; // -258
storage[3149] = -12'b000010101100; // -172
storage[3150] =  12'b000010001001; // 137
storage[3151] = -12'b000001010000; // -80
storage[3152] = -12'b000011011001; // -217
storage[3153] = -12'b000100011101; // -285
storage[3154] = -12'b000010010001; // -145
storage[3155] = -12'b000000011010; // -26
storage[3156] =  12'b000001001100; // 76
storage[3157] = -12'b000000111110; // -62
storage[3158] = -12'b000000011100; // -28
storage[3159] = -12'b000001001111; // -79
storage[3160] = -12'b000100011100; // -284
storage[3161] = -12'b000100101111; // -303
storage[3162] = -12'b000010100000; // -160
storage[3163] = -12'b001001010101; // -597
storage[3164] = -12'b000001000010; // -66
storage[3165] = -12'b000010100010; // -162
storage[3166] =  12'b000000011000; // 24
storage[3167] = -12'b000010010011; // -147
storage[3168] =  12'b000000011010; // 26
storage[3169] =  12'b000000001110; // 14
storage[3170] =  12'b000001001101; // 77
storage[3171] =  12'b000001011011; // 91
storage[3172] =  12'b000011111011; // 251
storage[3173] =  12'b000001110101; // 117
storage[3174] =  12'b000000000001; // 1
storage[3175] =  12'b000001101110; // 110
storage[3176] =  12'b000001101000; // 104
storage[3177] = -12'b000100000000; // -256
storage[3178] = -12'b000011101101; // -237
storage[3179] = -12'b000100101100; // -300
storage[3180] =  12'b000000101000; // 40
storage[3181] =  12'b000010011001; // 153
storage[3182] = -12'b000001001111; // -79
storage[3183] =  12'b000000111100; // 60
storage[3184] = -12'b000001111011; // -123
storage[3185] = -12'b000010100100; // -164
storage[3186] = -12'b000010101000; // -168
storage[3187] = -12'b000110111110; // -446
storage[3188] = -12'b000111111110; // -510
storage[3189] = -12'b000100111000; // -312
storage[3190] =  12'b000100100110; // 294
storage[3191] =  12'b000010111110; // 190
storage[3192] = -12'b000000000110; // -6
storage[3193] = -12'b000100001111; // -271
storage[3194] = -12'b000000110101; // -53
storage[3195] = -12'b000000010100; // -20
storage[3196] = -12'b001000100101; // -549
storage[3197] = -12'b000111111101; // -509
storage[3198] = -12'b000010001101; // -141
storage[3199] =  12'b000001001100; // 76
storage[3200] = -12'b000010100101; // -165
storage[3201] = -12'b000011010111; // -215
storage[3202] =  12'b000010100101; // 165
storage[3203] = -12'b000000100010; // -34
storage[3204] = -12'b000011011001; // -217
storage[3205] =  12'b000000101100; // 44
storage[3206] = -12'b000010001100; // -140
storage[3207] =  12'b000010010011; // 147
storage[3208] = -12'b000001000100; // -68
storage[3209] =  12'b000001100101; // 101
storage[3210] = -12'b000000011001; // -25
storage[3211] =  12'b000000101100; // 44
storage[3212] = -12'b000000100001; // -33
storage[3213] = -12'b001000000011; // -515
storage[3214] = -12'b000001111001; // -121
storage[3215] = -12'b000100101010; // -298
storage[3216] = -12'b000100001000; // -264
storage[3217] = -12'b000000111100; // -60
storage[3218] = -12'b000001000010; // -66
storage[3219] = -12'b000010011000; // -152
storage[3220] = -12'b000000111011; // -59
storage[3221] =  12'b000001001111; // 79
storage[3222] =  12'b000001000001; // 65
storage[3223] = -12'b000111001101; // -461
storage[3224] = -12'b000100011111; // -287
storage[3225] = -12'b000000111100; // -60
storage[3226] = -12'b000000011100; // -28
storage[3227] = -12'b000001100111; // -103
storage[3228] = -12'b000001010101; // -85
storage[3229] =  12'b000010001000; // 136
storage[3230] = -12'b000001010101; // -85
storage[3231] = -12'b000000101011; // -43
storage[3232] = -12'b000001111101; // -125
storage[3233] = -12'b000010001001; // -137
storage[3234] = -12'b000001010100; // -84
storage[3235] = -12'b000010100100; // -164
storage[3236] = -12'b000001100111; // -103
storage[3237] = -12'b000000101011; // -43
storage[3238] = -12'b000010011010; // -154
storage[3239] = -12'b000000011000; // -24
storage[3240] = -12'b000000101010; // -42
storage[3241] =  12'b000000110101; // 53
storage[3242] = -12'b000010001110; // -142
storage[3243] =  12'b000001110011; // 115
storage[3244] = -12'b000100001001; // -265
storage[3245] = -12'b000010001000; // -136
storage[3246] =  12'b000000011001; // 25
storage[3247] = -12'b000110001011; // -395
storage[3248] =  12'b000010010101; // 149
storage[3249] =  12'b000010110000; // 176
storage[3250] = -12'b000001111001; // -121
storage[3251] =  12'b000000010100; // 20
storage[3252] =  12'b000001010011; // 83
storage[3253] =  12'b000100000011; // 259
storage[3254] =  12'b000001011110; // 94
storage[3255] = -12'b000001110001; // -113
storage[3256] = -12'b000011010001; // -209
storage[3257] = -12'b000011011110; // -222
storage[3258] = -12'b000000110001; // -49
storage[3259] =  12'b000001010001; // 81
storage[3260] = -12'b000000010010; // -18
storage[3261] =  12'b000011000001; // 193
storage[3262] =  12'b000100000110; // 262
storage[3263] = -12'b000001011000; // -88
storage[3264] =  12'b000000100001; // 33
storage[3265] =  12'b000001010010; // 82
storage[3266] = -12'b000001100000; // -96
storage[3267] = -12'b000110000110; // -390
storage[3268] = -12'b000001001001; // -73
storage[3269] = -12'b000001101010; // -106
storage[3270] = -12'b000001010011; // -83
storage[3271] =  12'b000000100101; // 37
storage[3272] =  12'b000000110111; // 55
storage[3273] = -12'b000010001000; // -136
storage[3274] = -12'b000000010001; // -17
storage[3275] = -12'b000000101010; // -42
storage[3276] =  12'b000000000001; // 1
storage[3277] = -12'b000000100101; // -37
storage[3278] = -12'b000010111001; // -185
storage[3279] = -12'b000010001000; // -136
storage[3280] = -12'b000000011111; // -31
storage[3281] = -12'b000010000100; // -132
storage[3282] =  12'b000000111011; // 59
storage[3283] = -12'b000001001100; // -76
storage[3284] = -12'b000011000010; // -194
storage[3285] =  12'b000000101110; // 46
storage[3286] =  12'b000000101000; // 40
storage[3287] = -12'b000001100110; // -102
storage[3288] = -12'b000000101110; // -46
storage[3289] = -12'b000000010000; // -16
storage[3290] = -12'b000000101100; // -44
storage[3291] =  12'b000001001101; // 77
storage[3292] = -12'b000000110001; // -49
storage[3293] = -12'b000010000100; // -132
storage[3294] =  12'b000000100110; // 38
storage[3295] =  12'b000000000100; // 4
storage[3296] =  12'b000000001000; // 8
storage[3297] = -12'b000010010011; // -147
storage[3298] = -12'b000000101100; // -44
storage[3299] =  12'b000000100011; // 35
storage[3300] = -12'b000000101001; // -41
storage[3301] =  12'b000001000111; // 71
storage[3302] = -12'b000000011111; // -31
storage[3303] = -12'b000010101111; // -175
storage[3304] =  12'b000000110010; // 50
storage[3305] =  12'b000000101001; // 41
storage[3306] =  12'b000000101001; // 41
storage[3307] = -12'b000001010011; // -83
storage[3308] = -12'b000001011001; // -89
storage[3309] =  12'b000000100001; // 33
storage[3310] = -12'b000001010111; // -87
storage[3311] = -12'b000011101001; // -233
storage[3312] = -12'b000010101000; // -168
storage[3313] = -12'b000001000010; // -66
storage[3314] = -12'b000010100100; // -164
storage[3315] = -12'b000010110010; // -178
storage[3316] =  12'b000000101011; // 43
storage[3317] = -12'b000011110101; // -245
storage[3318] = -12'b000010000001; // -129
storage[3319] = -12'b000000010001; // -17
storage[3320] = -12'b000011001001; // -201
storage[3321] =  12'b000000111010; // 58
storage[3322] =  12'b000000101001; // 41
storage[3323] = -12'b000011000000; // -192
storage[3324] =  12'b000001001011; // 75
storage[3325] =  12'b000001101011; // 107
storage[3326] = -12'b000001111100; // -124
storage[3327] = -12'b000000000100; // -4
storage[3328] = -12'b000010011001; // -153
storage[3329] =  12'b000000001110; // 14
storage[3330] =  12'b000000010000; // 16
storage[3331] = -12'b000000011101; // -29
storage[3332] = -12'b000001001110; // -78
storage[3333] = -12'b000000001100; // -12
storage[3334] = -12'b000010000011; // -131
storage[3335] = -12'b000001011000; // -88
storage[3336] =  12'b000001001010; // 74
storage[3337] = -12'b000000011000; // -24
storage[3338] =  12'b000001011000; // 88
storage[3339] = -12'b000010010111; // -151
storage[3340] = -12'b000001110001; // -113
storage[3341] =  12'b000000101110; // 46
storage[3342] =  12'b000000000010; // 2
storage[3343] =  12'b000000011011; // 27
storage[3344] =  12'b000000011111; // 31
storage[3345] = -12'b000011101011; // -235
storage[3346] =  12'b000000110010; // 50
storage[3347] =  12'b000000001010; // 10
storage[3348] =  12'b000000101011; // 43
storage[3349] = -12'b000010101101; // -173
storage[3350] = -12'b000010101101; // -173
storage[3351] = -12'b000001010111; // -87
storage[3352] = -12'b000010011111; // -159
storage[3353] = -12'b000000110101; // -53
storage[3354] =  12'b000001011010; // 90
storage[3355] = -12'b000010011111; // -159
storage[3356] = -12'b000001000010; // -66
storage[3357] = -12'b000001110110; // -118
storage[3358] = -12'b000000010000; // -16
storage[3359] =  12'b000000111101; // 61
storage[3360] =  12'b000001000000; // 64
storage[3361] = -12'b000010010010; // -146
storage[3362] =  12'b000000110110; // 54
storage[3363] = -12'b000000011011; // -27
storage[3364] = -12'b000010001110; // -142
storage[3365] = -12'b000001101010; // -106
storage[3366] =  12'b000000111111; // 63
storage[3367] = -12'b000000010001; // -17
storage[3368] =  12'b000000011110; // 30
storage[3369] = -12'b000000101011; // -43
storage[3370] = -12'b000001010010; // -82
storage[3371] =  12'b000000010111; // 23
storage[3372] = -12'b000010010011; // -147
storage[3373] = -12'b000001010010; // -82
storage[3374] = -12'b000010100010; // -162
storage[3375] = -12'b000000111110; // -62
storage[3376] = -12'b000000001001; // -9
storage[3377] = -12'b000000111000; // -56
storage[3378] = -12'b000010110011; // -179
storage[3379] = -12'b000001001001; // -73
storage[3380] = -12'b000011000000; // -192
storage[3381] = -12'b000001110100; // -116
storage[3382] = -12'b000010011111; // -159
storage[3383] = -12'b000001100110; // -102
storage[3384] =  12'b000000101010; // 42
storage[3385] =  12'b000000110101; // 53
storage[3386] = -12'b000001000111; // -71
storage[3387] = -12'b000000110010; // -50
storage[3388] = -12'b000010110110; // -182
storage[3389] =  12'b000000001101; // 13
storage[3390] = -12'b000001101101; // -109
storage[3391] =  12'b000000000110; // 6
storage[3392] =  12'b000001010101; // 85
storage[3393] = -12'b000001001110; // -78
storage[3394] = -12'b000001110100; // -116
storage[3395] = -12'b000001110101; // -117
storage[3396] =  12'b000000001110; // 14
storage[3397] =  12'b000001000011; // 67
storage[3398] =  12'b000000100100; // 36
storage[3399] = -12'b000001010011; // -83
storage[3400] =  12'b000001110001; // 113
storage[3401] =  12'b000000010110; // 22
storage[3402] =  12'b000001100000; // 96
storage[3403] = -12'b000000011100; // -28
storage[3404] = -12'b000000100011; // -35
storage[3405] = -12'b000010000110; // -134
storage[3406] =  12'b000000000011; // 3
storage[3407] = -12'b000000000110; // -6
storage[3408] = -12'b000000001010; // -10
storage[3409] = -12'b000001100100; // -100
storage[3410] = -12'b000001011111; // -95
storage[3411] =  12'b000000011111; // 31
storage[3412] =  12'b000000011100; // 28
storage[3413] = -12'b000000100101; // -37
storage[3414] =  12'b000000001000; // 8
storage[3415] =  12'b000010100001; // 161
storage[3416] =  12'b000000010110; // 22
storage[3417] =  12'b000000110111; // 55
storage[3418] = -12'b001000010011; // -531
storage[3419] =  12'b000000001010; // 10
storage[3420] =  12'b000011010010; // 210
storage[3421] =  12'b000010101101; // 173
storage[3422] =  12'b000001110001; // 113
storage[3423] =  12'b000001100011; // 99
storage[3424] =  12'b000011000011; // 195
storage[3425] =  12'b000010000010; // 130
storage[3426] = -12'b000001010010; // -82
storage[3427] =  12'b000001111110; // 126
storage[3428] =  12'b000001111000; // 120
storage[3429] = -12'b000001111000; // -120
storage[3430] = -12'b001000110101; // -565
storage[3431] = -12'b001001110100; // -628
storage[3432] = -12'b000010111111; // -191
storage[3433] =  12'b000011110001; // 241
storage[3434] = -12'b000000000110; // -6
storage[3435] = -12'b000001111100; // -124
storage[3436] = -12'b000111011000; // -472
storage[3437] = -12'b000011011000; // -216
storage[3438] =  12'b000001011010; // 90
storage[3439] =  12'b000000111101; // 61
storage[3440] = -12'b000010001001; // -137
storage[3441] = -12'b000110110110; // -438
storage[3442] =  12'b000010001110; // 142
storage[3443] =  12'b000000000100; // 4
storage[3444] =  12'b000000111100; // 60
storage[3445] = -12'b000011000000; // -192
storage[3446] =  12'b000100001101; // 269
storage[3447] =  12'b000001001010; // 74
storage[3448] = -12'b000010011000; // -152
storage[3449] = -12'b000010100001; // -161
storage[3450] =  12'b000000110011; // 51
storage[3451] =  12'b000000010001; // 17
storage[3452] =  12'b000011111010; // 250
storage[3453] =  12'b000000011110; // 30
storage[3454] = -12'b000001011110; // -94
storage[3455] = -12'b000001100000; // -96
storage[3456] = -12'b000010000000; // -128
storage[3457] = -12'b000011101100; // -236
storage[3458] = -12'b000010000000; // -128
storage[3459] = -12'b000000000100; // -4
storage[3460] =  12'b000011000100; // 196
storage[3461] = -12'b000000011110; // -30
storage[3462] = -12'b000011001100; // -204
storage[3463] =  12'b000001000110; // 70
storage[3464] = -12'b000000001010; // -10
storage[3465] = -12'b000110010011; // -403
storage[3466] =  12'b000010111010; // 186
storage[3467] =  12'b000000111010; // 58
storage[3468] = -12'b000001101111; // -111
storage[3469] = -12'b000000011111; // -31
storage[3470] = -12'b000000010000; // -16
storage[3471] =  12'b000000000001; // 1
storage[3472] =  12'b000000101111; // 47
storage[3473] = -12'b000010011001; // -153
storage[3474] = -12'b000011001010; // -202
storage[3475] = -12'b001011010111; // -727
storage[3476] = -12'b000110110010; // -434
storage[3477] = -12'b000111000101; // -453
storage[3478] =  12'b000010011001; // 153
storage[3479] =  12'b000101001000; // 328
storage[3480] = -12'b000100110100; // -308
storage[3481] = -12'b000001000100; // -68
storage[3482] = -12'b000010001111; // -143
storage[3483] = -12'b000000001111; // -15
storage[3484] = -12'b000100001110; // -270
storage[3485] = -12'b000110011001; // -409
storage[3486] = -12'b001001100110; // -614
storage[3487] = -12'b000000001110; // -14
storage[3488] = -12'b000000001111; // -15
storage[3489] = -12'b001001001100; // -588
storage[3490] =  12'b000011011001; // 217
storage[3491] =  12'b000010110111; // 183
storage[3492] =  12'b000001001001; // 73
storage[3493] =  12'b000011011111; // 223
storage[3494] =  12'b000001100001; // 97
storage[3495] = -12'b000000100101; // -37
storage[3496] = -12'b000001010101; // -85
storage[3497] =  12'b000000100000; // 32
storage[3498] = -12'b000010100011; // -163
storage[3499] = -12'b000000100111; // -39
storage[3500] =  12'b000000101010; // 42
storage[3501] = -12'b000010101111; // -175
storage[3502] =  12'b000010000011; // 131
storage[3503] = -12'b000011010011; // -211
storage[3504] = -12'b000100100010; // -290
storage[3505] =  12'b000000100101; // 37
storage[3506] =  12'b000011001110; // 206
storage[3507] = -12'b000001000001; // -65
storage[3508] =  12'b000010110010; // 178
storage[3509] =  12'b000001010110; // 86
storage[3510] =  12'b000001011011; // 91
storage[3511] = -12'b000011011000; // -216
storage[3512] =  12'b000001010110; // 86
storage[3513] = -12'b000011010000; // -208
storage[3514] = -12'b000000010010; // -18
storage[3515] = -12'b000000100011; // -35
storage[3516] = -12'b000000001100; // -12
storage[3517] =  12'b000000001011; // 11
storage[3518] =  12'b000001010000; // 80
storage[3519] =  12'b000000001010; // 10
storage[3520] = -12'b000011001110; // -206
storage[3521] = -12'b000101010010; // -338
storage[3522] = -12'b000001110010; // -114
storage[3523] =  12'b000001111100; // 124
storage[3524] = -12'b000010010001; // -145
storage[3525] = -12'b000000101000; // -40
storage[3526] =  12'b000000111101; // 61
storage[3527] =  12'b000010011010; // 154
storage[3528] = -12'b000101011100; // -348
storage[3529] = -12'b000001000110; // -70
storage[3530] =  12'b000000110100; // 52
storage[3531] =  12'b000000101000; // 40
storage[3532] = -12'b000111000010; // -450
storage[3533] =  12'b000000000100; // 4
storage[3534] =  12'b000001101011; // 107
storage[3535] = -12'b000010001010; // -138
storage[3536] =  12'b000010110100; // 180
storage[3537] =  12'b000010110000; // 176
storage[3538] = -12'b000100000101; // -261
storage[3539] =  12'b000001100011; // 99
storage[3540] =  12'b000000001100; // 12
storage[3541] = -12'b000001010101; // -85
storage[3542] = -12'b000000010011; // -19
storage[3543] = -12'b000011111000; // -248
storage[3544] =  12'b000000111111; // 63
storage[3545] = -12'b000001100010; // -98
storage[3546] =  12'b000001001111; // 79
storage[3547] = -12'b000000110011; // -51
storage[3548] = -12'b000000101000; // -40
storage[3549] = -12'b000000110011; // -51
storage[3550] =  12'b000001101110; // 110
storage[3551] =  12'b000001000111; // 71
storage[3552] = -12'b000011011011; // -219
storage[3553] =  12'b000010000001; // 129
storage[3554] =  12'b000000110000; // 48
storage[3555] = -12'b000100010011; // -275
storage[3556] = -12'b000000110001; // -49
storage[3557] =  12'b000000011001; // 25
storage[3558] = -12'b000100001011; // -267
storage[3559] =  12'b000000111111; // 63
storage[3560] = -12'b000101100011; // -355
storage[3561] = -12'b000101000110; // -326
storage[3562] = -12'b000000000100; // -4
storage[3563] =  12'b000000001011; // 11
storage[3564] =  12'b000100001011; // 267
storage[3565] =  12'b000001000010; // 66
storage[3566] =  12'b000000001011; // 11
storage[3567] = -12'b000000101000; // -40
storage[3568] =  12'b000100000010; // 258
storage[3569] =  12'b000010001010; // 138
storage[3570] = -12'b000000010011; // -19
storage[3571] =  12'b000001000111; // 71
storage[3572] =  12'b000001100010; // 98
storage[3573] =  12'b000001111111; // 127
storage[3574] = -12'b000000000100; // -4
storage[3575] =  12'b000010000110; // 134
storage[3576] = -12'b000001010110; // -86
storage[3577] = -12'b000010101100; // -172
storage[3578] = -12'b000001100010; // -98
storage[3579] = -12'b001011011010; // -730
storage[3580] = -12'b000000101100; // -44
storage[3581] = -12'b001010100101; // -677
storage[3582] =  12'b000011111100; // 252
storage[3583] =  12'b000010100111; // 167
storage[3584] =  12'b000001001011; // 75
storage[3585] =  12'b000001111010; // 122
storage[3586] = -12'b000001111000; // -120
storage[3587] =  12'b000010001110; // 142
storage[3588] =  12'b000000111101; // 61
storage[3589] = -12'b000011101110; // -238
storage[3590] = -12'b000000000100; // -4
storage[3591] =  12'b000000011100; // 28
storage[3592] =  12'b000011011110; // 222
storage[3593] =  12'b000010000101; // 133
storage[3594] = -12'b000010001100; // -140
storage[3595] =  12'b000000111001; // 57
storage[3596] = -12'b000001000010; // -66
storage[3597] =  12'b000010000010; // 130
storage[3598] = -12'b000000110101; // -53
storage[3599] = -12'b000110011001; // -409
storage[3600] = -12'b000000111101; // -61
storage[3601] = -12'b000011010110; // -214
storage[3602] =  12'b000010001010; // 138
storage[3603] =  12'b000011010001; // 209
storage[3604] =  12'b000000101001; // 41
storage[3605] =  12'b000001111111; // 127
storage[3606] = -12'b000011011111; // -223
storage[3607] = -12'b000000001111; // -15
storage[3608] = -12'b000000011110; // -30
storage[3609] =  12'b000010101111; // 175
storage[3610] = -12'b000000100011; // -35
storage[3611] =  12'b000001100100; // 100
storage[3612] =  12'b000000101000; // 40
storage[3613] =  12'b000010100100; // 164
storage[3614] =  12'b000001000111; // 71
storage[3615] = -12'b000010011001; // -153
storage[3616] =  12'b000001010110; // 86
storage[3617] =  12'b000000110100; // 52
storage[3618] =  12'b000000100000; // 32
storage[3619] = -12'b000010010000; // -144
storage[3620] = -12'b000001110101; // -117
storage[3621] = -12'b000010100010; // -162
storage[3622] =  12'b000001011010; // 90
storage[3623] =  12'b000100101111; // 303
storage[3624] =  12'b000000011101; // 29
storage[3625] = -12'b000000010110; // -22
storage[3626] =  12'b000001000010; // 66
storage[3627] =  12'b000100000001; // 257
storage[3628] = -12'b000001000001; // -65
storage[3629] =  12'b000010010001; // 145
storage[3630] =  12'b000010111110; // 190
storage[3631] =  12'b000000010111; // 23
storage[3632] =  12'b000001111011; // 123
storage[3633] =  12'b000001100011; // 99
storage[3634] = -12'b000000101111; // -47
storage[3635] =  12'b000000000010; // 2
storage[3636] =  12'b000010000110; // 134
storage[3637] =  12'b000011001101; // 205
storage[3638] =  12'b000000101100; // 44
storage[3639] =  12'b000010001111; // 143
storage[3640] =  12'b000010100001; // 161
storage[3641] =  12'b000010000110; // 134
storage[3642] =  12'b000010000111; // 135
storage[3643] =  12'b000011001111; // 207
storage[3644] =  12'b000011001100; // 204
storage[3645] = -12'b000001010000; // -80
storage[3646] = -12'b000001000100; // -68
storage[3647] = -12'b000010010001; // -145
storage[3648] =  12'b000011110010; // 242
storage[3649] =  12'b000001011101; // 93
storage[3650] =  12'b000000011111; // 31
storage[3651] = -12'b000000000111; // -7
storage[3652] =  12'b000001111100; // 124
storage[3653] = -12'b000100111111; // -319
storage[3654] = -12'b000011101001; // -233
storage[3655] =  12'b000000001100; // 12
storage[3656] =  12'b000001101110; // 110
storage[3657] = -12'b000010010111; // -151
storage[3658] = -12'b000011110000; // -240
storage[3659] = -12'b000000111101; // -61
storage[3660] = -12'b000011001011; // -203
storage[3661] =  12'b000101100111; // 359
storage[3662] =  12'b000011111010; // 250
storage[3663] =  12'b000011011100; // 220
storage[3664] = -12'b000000000110; // -6
storage[3665] =  12'b000011110110; // 246
storage[3666] =  12'b000100100010; // 290
storage[3667] = -12'b000000011010; // -26
storage[3668] = -12'b000000101110; // -46
storage[3669] =  12'b000011010011; // 211
storage[3670] =  12'b000010001011; // 139
storage[3671] = -12'b000000001110; // -14
storage[3672] = -12'b000010101011; // -171
storage[3673] = -12'b000001110110; // -118
storage[3674] = -12'b000101111011; // -379
storage[3675] = -12'b000101001110; // -334
storage[3676] = -12'b001000010001; // -529
storage[3677] = -12'b000100100111; // -295
storage[3678] =  12'b000100110100; // 308
storage[3679] =  12'b000001101100; // 108
storage[3680] = -12'b000000001111; // -15
storage[3681] = -12'b000001011011; // -91
storage[3682] =  12'b000011001101; // 205
storage[3683] =  12'b000011011001; // 217
storage[3684] = -12'b000001000111; // -71
storage[3685] = -12'b000000100001; // -33
storage[3686] = -12'b001001000011; // -579
storage[3687] = -12'b000010101111; // -175
storage[3688] = -12'b000011010000; // -208
storage[3689] = -12'b001000111100; // -572
storage[3690] = -12'b000110111111; // -447
storage[3691] =  12'b000001001001; // 73
storage[3692] = -12'b000000100111; // -39
storage[3693] = -12'b000001110011; // -115
storage[3694] =  12'b000000001001; // 9
storage[3695] = -12'b000000011111; // -31
storage[3696] =  12'b000000001000; // 8
storage[3697] =  12'b000000000010; // 2
storage[3698] =  12'b000000101111; // 47
storage[3699] =  12'b000000111001; // 57
storage[3700] =  12'b000110100011; // 419
storage[3701] =  12'b000000010001; // 17
storage[3702] =  12'b000001011100; // 92
storage[3703] = -12'b000000011111; // -31
storage[3704] = -12'b000010110100; // -180
storage[3705] = -12'b000000001101; // -13
storage[3706] = -12'b000110101011; // -427
storage[3707] =  12'b000000110111; // 55
storage[3708] =  12'b000000000101; // 5
storage[3709] = -12'b000001010111; // -87
storage[3710] = -12'b000000011001; // -25
storage[3711] = -12'b000010110001; // -177
storage[3712] = -12'b000001110111; // -119
storage[3713] = -12'b000001010110; // -86
storage[3714] = -12'b000010101111; // -175
storage[3715] = -12'b000000001111; // -15
storage[3716] = -12'b000100100101; // -293
storage[3717] = -12'b001010110011; // -691
storage[3718] = -12'b000001001000; // -72
storage[3719] = -12'b000011100101; // -229
storage[3720] =  12'b000001101110; // 110
storage[3721] = -12'b000100011110; // -286
storage[3722] = -12'b000010001110; // -142
storage[3723] =  12'b000001101000; // 104
storage[3724] =  12'b000010001101; // 141
storage[3725] =  12'b000000010010; // 18
storage[3726] =  12'b000010101110; // 174
storage[3727] = -12'b000001001011; // -75
storage[3728] =  12'b000001001010; // 74
storage[3729] =  12'b000001000011; // 67
storage[3730] =  12'b000100110111; // 311
storage[3731] =  12'b000010011101; // 157
storage[3732] =  12'b000011110001; // 241
storage[3733] =  12'b000100000011; // 259
storage[3734] =  12'b000001110110; // 118
storage[3735] =  12'b000010000110; // 134
storage[3736] =  12'b000011101111; // 239
storage[3737] = -12'b000000010111; // -23
storage[3738] =  12'b000010100000; // 160
storage[3739] =  12'b000011000011; // 195
storage[3740] =  12'b000000101110; // 46
storage[3741] =  12'b000011010001; // 209
storage[3742] =  12'b000100110101; // 309
storage[3743] =  12'b000001100101; // 101
storage[3744] =  12'b000101110001; // 369
storage[3745] =  12'b000010010110; // 150
storage[3746] = -12'b000000010101; // -21
storage[3747] = -12'b000000100111; // -39
storage[3748] = -12'b000001100000; // -96
storage[3749] =  12'b000000110000; // 48
storage[3750] = -12'b000001100001; // -97
storage[3751] = -12'b000001010011; // -83
storage[3752] =  12'b000001110000; // 112
storage[3753] =  12'b000000011011; // 27
storage[3754] = -12'b000000110001; // -49
storage[3755] =  12'b000001101101; // 109
storage[3756] =  12'b000011011110; // 222
storage[3757] =  12'b000001010111; // 87
storage[3758] =  12'b000101010101; // 341
storage[3759] =  12'b000101010010; // 338
storage[3760] =  12'b000011010100; // 212
storage[3761] =  12'b000000101010; // 42
storage[3762] =  12'b000110111000; // 440
storage[3763] =  12'b000001011000; // 88
storage[3764] =  12'b000000100000; // 32
storage[3765] =  12'b000001000100; // 68
storage[3766] =  12'b000000011101; // 29
storage[3767] =  12'b000000101010; // 42
storage[3768] =  12'b000000000100; // 4
storage[3769] =  12'b000001001010; // 74
storage[3770] =  12'b000010110011; // 179
storage[3771] =  12'b000000001101; // 13
storage[3772] =  12'b000100101101; // 301
storage[3773] =  12'b000011010111; // 215
storage[3774] =  12'b000010000101; // 133
storage[3775] =  12'b000010011100; // 156
storage[3776] = -12'b000000000111; // -7
storage[3777] = -12'b000011010111; // -215
storage[3778] = -12'b000011001111; // -207
storage[3779] = -12'b000011010011; // -211
storage[3780] = -12'b000010110110; // -182
storage[3781] = -12'b000001000101; // -69
storage[3782] =  12'b000000110000; // 48
storage[3783] =  12'b000001110101; // 117
storage[3784] =  12'b000000101011; // 43
storage[3785] =  12'b000001000000; // 64
storage[3786] =  12'b000101011000; // 344
storage[3787] = -12'b000010110000; // -176
storage[3788] =  12'b000000000011; // 3
storage[3789] =  12'b000010101111; // 175
storage[3790] = -12'b000000001010; // -10
storage[3791] =  12'b000000001001; // 9
storage[3792] =  12'b000001000010; // 66
storage[3793] =  12'b000100101101; // 301
storage[3794] =  12'b000000000010; // 2
storage[3795] = -12'b000000010101; // -21
storage[3796] = -12'b000010101101; // -173
storage[3797] = -12'b000011011101; // -221
storage[3798] = -12'b000000011000; // -24
storage[3799] = -12'b000001111110; // -126
storage[3800] = -12'b000001010100; // -84
storage[3801] = -12'b000000101100; // -44
storage[3802] =  12'b000101110011; // 371
storage[3803] =  12'b000001110101; // 117
storage[3804] = -12'b000000001111; // -15
storage[3805] = -12'b000010101000; // -168
storage[3806] =  12'b000000000001; // 1
storage[3807] = -12'b000000011011; // -27
storage[3808] =  12'b000000100000; // 32
storage[3809] = -12'b000101001101; // -333
storage[3810] = -12'b000000101000; // -40
storage[3811] =  12'b000001011011; // 91
storage[3812] = -12'b000111100001; // -481
storage[3813] =  12'b000001000100; // 68
storage[3814] =  12'b000000000000; // 0
storage[3815] = -12'b000011011100; // -220
storage[3816] = -12'b000000110011; // -51
storage[3817] =  12'b000011110110; // 246
storage[3818] =  12'b000010110110; // 182
storage[3819] =  12'b000010110111; // 183
storage[3820] =  12'b000001011001; // 89
storage[3821] =  12'b000000011100; // 28
storage[3822] =  12'b000000011111; // 31
storage[3823] = -12'b000011110110; // -246
storage[3824] = -12'b000011001101; // -205
storage[3825] =  12'b000000000010; // 2
storage[3826] = -12'b000011000001; // -193
storage[3827] = -12'b000000101111; // -47
storage[3828] =  12'b000011100000; // 224
storage[3829] =  12'b000001110011; // 115
storage[3830] =  12'b000010000101; // 133
storage[3831] =  12'b000100101101; // 301
storage[3832] =  12'b000001110110; // 118
storage[3833] = -12'b000000100101; // -37
storage[3834] =  12'b000010111111; // 191
storage[3835] =  12'b000100010100; // 276
storage[3836] =  12'b000100011100; // 284
storage[3837] =  12'b000101000011; // 323
storage[3838] =  12'b000000000101; // 5
storage[3839] =  12'b000000101000; // 40
storage[3840] = -12'b000101011001; // -345
storage[3841] = -12'b000100000101; // -261
storage[3842] = -12'b000110111001; // -441
storage[3843] = -12'b000111000000; // -448
storage[3844] = -12'b000001001001; // -73
storage[3845] = -12'b000000111010; // -58
storage[3846] =  12'b000000011101; // 29
storage[3847] = -12'b000001011011; // -91
storage[3848] = -12'b000000011110; // -30
storage[3849] =  12'b000011010110; // 214
storage[3850] =  12'b000100010101; // 277
storage[3851] =  12'b000100101111; // 303
storage[3852] = -12'b000000100010; // -34
storage[3853] = -12'b000000100011; // -35
storage[3854] =  12'b000001100110; // 102
storage[3855] =  12'b000010110101; // 181
storage[3856] = -12'b000100001001; // -265
storage[3857] = -12'b000101111110; // -382
storage[3858] =  12'b000011000000; // 192
storage[3859] = -12'b000101000110; // -326
storage[3860] =  12'b000000110011; // 51
storage[3861] =  12'b000000010010; // 18
storage[3862] = -12'b000000000010; // -2
storage[3863] = -12'b000000101111; // -47
storage[3864] = -12'b000000001111; // -15
storage[3865] = -12'b000010010001; // -145
storage[3866] = -12'b000010011011; // -155
storage[3867] =  12'b000000100100; // 36
storage[3868] =  12'b000010010101; // 149
storage[3869] =  12'b000000010000; // 16
storage[3870] = -12'b000001100011; // -99
storage[3871] = -12'b000001100000; // -96
storage[3872] =  12'b000000100111; // 39
storage[3873] =  12'b000001101001; // 105
storage[3874] = -12'b000001011110; // -94
storage[3875] =  12'b000001001000; // 72
storage[3876] = -12'b000001000101; // -69
storage[3877] =  12'b000100110100; // 308
storage[3878] =  12'b000010110100; // 180
storage[3879] = -12'b000010000000; // -128
storage[3880] =  12'b000011110111; // 247
storage[3881] =  12'b000011000001; // 193
storage[3882] =  12'b000010000001; // 129
storage[3883] = -12'b000010110011; // -179
storage[3884] = -12'b000001001010; // -74
storage[3885] = -12'b000010001111; // -143
storage[3886] = -12'b000101010001; // -337
storage[3887] = -12'b000000101010; // -42
storage[3888] =  12'b000010101111; // 175
storage[3889] =  12'b000000001011; // 11
storage[3890] =  12'b000000010110; // 22
storage[3891] = -12'b000010001011; // -139
storage[3892] = -12'b000000110001; // -49
storage[3893] = -12'b000000010111; // -23
storage[3894] = -12'b000010100110; // -166
storage[3895] =  12'b000000001010; // 10
storage[3896] = -12'b000000001001; // -9
storage[3897] =  12'b000001111110; // 126
storage[3898] =  12'b000010011111; // 159
storage[3899] =  12'b000010000011; // 131
storage[3900] = -12'b000000011101; // -29
storage[3901] =  12'b000001101000; // 104
storage[3902] =  12'b000011001011; // 203
storage[3903] =  12'b000000110001; // 49
storage[3904] =  12'b000000010100; // 20
storage[3905] = -12'b000000001001; // -9
storage[3906] =  12'b000111101010; // 490
storage[3907] =  12'b000001001100; // 76
storage[3908] = -12'b000000111100; // -60
storage[3909] = -12'b000011011000; // -216
storage[3910] =  12'b000001000100; // 68
storage[3911] =  12'b000001101101; // 109
storage[3912] = -12'b000011101101; // -237
storage[3913] = -12'b000000011101; // -29
storage[3914] = -12'b000000001001; // -9
storage[3915] =  12'b000000000111; // 7
storage[3916] = -12'b000010000000; // -128
storage[3917] = -12'b000001101011; // -107
storage[3918] = -12'b000011101111; // -239
storage[3919] =  12'b000100000010; // 258
storage[3920] = -12'b000000000011; // -3
storage[3921] = -12'b000010011001; // -153
storage[3922] =  12'b000101011011; // 347
storage[3923] =  12'b000100011011; // 283
storage[3924] =  12'b000001011111; // 95
storage[3925] =  12'b000010110001; // 177
storage[3926] = -12'b000010011111; // -159
storage[3927] = -12'b000011010000; // -208
storage[3928] =  12'b000000111010; // 58
storage[3929] = -12'b000010110100; // -180
storage[3930] = -12'b000010100000; // -160
storage[3931] = -12'b000101110001; // -369
storage[3932] = -12'b001111111101; // -1021
storage[3933] = -12'b000000010101; // -21
storage[3934] =  12'b000010010110; // 150
storage[3935] = -12'b000000101101; // -45
storage[3936] = -12'b000001011110; // -94
storage[3937] =  12'b000001001101; // 77
storage[3938] = -12'b000000100101; // -37
storage[3939] = -12'b000011000000; // -192
storage[3940] = -12'b000101100110; // -358
storage[3941] = -12'b000111110101; // -501
storage[3942] = -12'b000001011111; // -95
storage[3943] =  12'b000001011110; // 94
storage[3944] =  12'b000001011111; // 95
storage[3945] =  12'b000001011000; // 88
storage[3946] =  12'b000000010010; // 18
storage[3947] = -12'b000001110110; // -118
storage[3948] =  12'b000001110110; // 118
storage[3949] = -12'b000001100010; // -98
storage[3950] = -12'b000000010101; // -21
storage[3951] =  12'b000010010100; // 148
storage[3952] =  12'b000101111110; // 382
storage[3953] = -12'b000010001100; // -140
storage[3954] = -12'b001000001111; // -527
storage[3955] =  12'b000011010011; // 211
storage[3956] = -12'b000010000001; // -129
storage[3957] = -12'b000010100011; // -163
storage[3958] =  12'b000001100001; // 97
storage[3959] = -12'b000001100100; // -100
storage[3960] = -12'b000010010000; // -144
storage[3961] =  12'b000010000010; // 130
storage[3962] =  12'b000000010010; // 18
storage[3963] = -12'b000000001111; // -15
storage[3964] = -12'b000000010111; // -23
storage[3965] =  12'b000000000000; // 0
storage[3966] =  12'b000000100001; // 33
storage[3967] =  12'b000001001111; // 79
storage[3968] = -12'b000011010000; // -208
storage[3969] = -12'b000000000111; // -7
storage[3970] =  12'b000011000100; // 196
storage[3971] =  12'b000100001110; // 270
storage[3972] =  12'b000011001010; // 202
storage[3973] =  12'b000000000011; // 3
storage[3974] =  12'b000011111010; // 250
storage[3975] =  12'b000000101010; // 42
storage[3976] =  12'b000011010010; // 210
storage[3977] =  12'b000010010110; // 150
storage[3978] = -12'b000000110101; // -53
storage[3979] = -12'b000001011101; // -93
storage[3980] = -12'b000000100110; // -38
storage[3981] = -12'b000001110111; // -119
storage[3982] = -12'b000001010010; // -82
storage[3983] = -12'b000011010100; // -212
storage[3984] =  12'b000001100100; // 100
storage[3985] =  12'b000010010110; // 150
storage[3986] = -12'b000001011111; // -95
storage[3987] =  12'b000000001101; // 13
storage[3988] = -12'b000000010101; // -21
storage[3989] =  12'b000000101100; // 44
storage[3990] = -12'b000010101000; // -168
storage[3991] = -12'b000001000001; // -65
storage[3992] = -12'b000000100001; // -33
storage[3993] =  12'b000001011000; // 88
storage[3994] = -12'b000000101000; // -40
storage[3995] =  12'b000000111100; // 60
storage[3996] =  12'b000010111111; // 191
storage[3997] = -12'b000011111011; // -251
storage[3998] = -12'b000010101001; // -169
storage[3999] =  12'b000001111001; // 121
storage[4000] = -12'b000011000110; // -198
storage[4001] =  12'b000010110011; // 179
storage[4002] =  12'b000001101111; // 111
storage[4003] = -12'b000001010111; // -87
storage[4004] =  12'b000100111011; // 315
storage[4005] =  12'b000100100111; // 295
storage[4006] =  12'b000000011100; // 28
storage[4007] =  12'b000010100111; // 167
storage[4008] =  12'b000010100100; // 164
storage[4009] =  12'b000001000010; // 66
storage[4010] =  12'b000001110100; // 116
storage[4011] = -12'b000000011110; // -30
storage[4012] =  12'b000001111111; // 127
storage[4013] = -12'b000011101011; // -235
storage[4014] =  12'b000100100111; // 295
storage[4015] =  12'b000011110000; // 240
storage[4016] = -12'b000001010001; // -81
storage[4017] = -12'b000000011101; // -29
storage[4018] =  12'b000010101001; // 169
storage[4019] =  12'b000001111100; // 124
storage[4020] =  12'b000100111010; // 314
storage[4021] = -12'b000100000000; // -256
storage[4022] =  12'b000110000101; // 389
storage[4023] =  12'b000010110101; // 181
storage[4024] =  12'b000001000110; // 70
storage[4025] = -12'b000000101011; // -43
storage[4026] = -12'b000000101100; // -44
storage[4027] =  12'b000001010100; // 84
storage[4028] = -12'b000011110101; // -245
storage[4029] = -12'b000100100011; // -291
storage[4030] =  12'b000010110111; // 183
storage[4031] = -12'b000010001011; // -139
storage[4032] =  12'b000000010101; // 21
storage[4033] =  12'b000000001011; // 11
storage[4034] = -12'b000000101001; // -41
storage[4035] =  12'b000000011000; // 24
storage[4036] = -12'b000000010000; // -16
storage[4037] =  12'b000000100101; // 37
storage[4038] = -12'b000010010010; // -146
storage[4039] = -12'b000000001100; // -12
storage[4040] = -12'b000011111001; // -249
storage[4041] = -12'b000011010100; // -212
storage[4042] = -12'b000010101000; // -168
storage[4043] = -12'b000000101111; // -47
storage[4044] = -12'b000001101100; // -108
storage[4045] = -12'b000010001000; // -136
storage[4046] =  12'b000001111110; // 126
storage[4047] =  12'b000010011011; // 155
storage[4048] =  12'b000000111101; // 61
storage[4049] =  12'b000000000110; // 6
storage[4050] =  12'b000000101110; // 46
storage[4051] = -12'b000000011010; // -26
storage[4052] =  12'b000001011101; // 93
storage[4053] = -12'b000100001101; // -269
storage[4054] =  12'b000000011100; // 28
storage[4055] = -12'b000001110110; // -118
storage[4056] = -12'b000011001110; // -206
storage[4057] = -12'b000010100100; // -164
storage[4058] = -12'b000000011011; // -27
storage[4059] =  12'b000000111001; // 57
storage[4060] =  12'b000010001010; // 138
storage[4061] = -12'b000010100001; // -161
storage[4062] =  12'b000000101110; // 46
storage[4063] = -12'b000001001011; // -75
storage[4064] = -12'b000000111010; // -58
storage[4065] = -12'b000001110101; // -117
storage[4066] = -12'b000010000001; // -129
storage[4067] =  12'b000011001111; // 207
storage[4068] = -12'b000000010001; // -17
storage[4069] =  12'b000010101100; // 172
storage[4070] = -12'b000011100111; // -231
storage[4071] =  12'b000000010111; // 23
storage[4072] =  12'b000000100000; // 32
storage[4073] =  12'b000001110001; // 113
storage[4074] =  12'b000001101011; // 107
storage[4075] =  12'b000010100101; // 165
storage[4076] =  12'b000100010001; // 273
storage[4077] =  12'b000010000011; // 131
storage[4078] = -12'b000001110010; // -114
storage[4079] = -12'b000100101101; // -301
storage[4080] = -12'b000000101010; // -42
storage[4081] =  12'b000000111101; // 61
storage[4082] =  12'b000000101111; // 47
storage[4083] =  12'b000110000010; // 386
storage[4084] =  12'b000000101100; // 44
storage[4085] =  12'b000001111100; // 124
storage[4086] =  12'b000011001011; // 203
storage[4087] =  12'b000000011100; // 28
storage[4088] = -12'b000010100011; // -163
storage[4089] = -12'b000101000100; // -324
storage[4090] =  12'b000000101101; // 45
storage[4091] = -12'b000000001000; // -8
storage[4092] =  12'b000000100010; // 34
storage[4093] =  12'b000010011100; // 156
storage[4094] = -12'b000000111101; // -61
storage[4095] =  12'b000011101011; // 235
storage[4096] = -12'b000010100110; // -166
storage[4097] = -12'b000001000100; // -68
storage[4098] = -12'b000001010101; // -85
storage[4099] = -12'b000011111010; // -250
storage[4100] = -12'b000001000101; // -69
storage[4101] =  12'b000001010001; // 81
storage[4102] = -12'b000000110101; // -53
storage[4103] =  12'b000000101000; // 40
storage[4104] =  12'b000000111011; // 59
storage[4105] =  12'b000010100100; // 164
storage[4106] =  12'b000001111101; // 125
storage[4107] =  12'b000001111110; // 126
storage[4108] = -12'b000001011101; // -93
storage[4109] = -12'b000000110111; // -55
storage[4110] =  12'b000001001101; // 77
storage[4111] = -12'b000001110111; // -119
storage[4112] = -12'b000010010110; // -150
storage[4113] =  12'b000001010010; // 82
storage[4114] = -12'b000001010100; // -84
storage[4115] =  12'b000001110111; // 119
storage[4116] =  12'b000100100100; // 292
storage[4117] = -12'b000010110011; // -179
storage[4118] = -12'b001110000100; // -900
storage[4119] = -12'b000011111000; // -248
storage[4120] =  12'b000010011100; // 156
storage[4121] = -12'b000100111000; // -312
storage[4122] = -12'b000001111101; // -125
storage[4123] =  12'b000001100010; // 98
storage[4124] = -12'b000001000110; // -70
storage[4125] = -12'b000011110001; // -241
storage[4126] = -12'b000011011111; // -223
storage[4127] = -12'b000011100111; // -231
storage[4128] =  12'b000000101010; // 42
storage[4129] = -12'b000001000111; // -71
storage[4130] =  12'b000000100110; // 38
storage[4131] =  12'b000010101100; // 172
storage[4132] = -12'b000001100001; // -97
storage[4133] =  12'b000001010011; // 83
storage[4134] =  12'b000011010001; // 209
storage[4135] = -12'b000100001100; // -268
storage[4136] =  12'b000000011010; // 26
storage[4137] = -12'b000101011110; // -350
storage[4138] =  12'b000101100101; // 357
storage[4139] =  12'b000000000011; // 3
storage[4140] = -12'b000010100010; // -162
storage[4141] =  12'b000001001011; // 75
storage[4142] = -12'b000000010100; // -20
storage[4143] = -12'b000010110010; // -178
storage[4144] =  12'b000010001001; // 137
storage[4145] =  12'b000010011011; // 155
storage[4146] = -12'b000000100000; // -32
storage[4147] =  12'b000101101010; // 362
storage[4148] =  12'b000010101100; // 172
storage[4149] =  12'b000100001111; // 271
storage[4150] = -12'b000010100110; // -166
storage[4151] =  12'b000010100001; // 161
storage[4152] =  12'b000011010100; // 212
storage[4153] =  12'b000001000100; // 68
storage[4154] =  12'b000010110100; // 180
storage[4155] =  12'b000101011110; // 350
storage[4156] = -12'b000011110001; // -241
storage[4157] = -12'b000010101100; // -172
storage[4158] = -12'b000001011100; // -92
storage[4159] = -12'b000001010110; // -86
storage[4160] =  12'b000011110110; // 246
storage[4161] = -12'b000011000110; // -198
storage[4162] = -12'b000110100111; // -423
storage[4163] = -12'b000011000100; // -196
storage[4164] = -12'b000000011111; // -31
storage[4165] = -12'b000100011101; // -285
storage[4166] = -12'b000010110110; // -182
storage[4167] = -12'b000000011001; // -25
storage[4168] =  12'b000010001111; // 143
storage[4169] =  12'b000000000100; // 4
storage[4170] =  12'b000000000111; // 7
storage[4171] =  12'b000011001100; // 204
storage[4172] = -12'b000001010111; // -87
storage[4173] =  12'b000101100101; // 357
storage[4174] = -12'b000000001101; // -13
storage[4175] = -12'b000000111001; // -57
storage[4176] = -12'b000010110011; // -179
storage[4177] = -12'b000001100110; // -102
storage[4178] = -12'b000000000010; // -2
storage[4179] =  12'b000000001010; // 10
storage[4180] =  12'b000001101000; // 104
storage[4181] =  12'b000010101100; // 172
storage[4182] =  12'b000011011101; // 221
storage[4183] =  12'b000000100011; // 35
storage[4184] =  12'b000010010001; // 145
storage[4185] =  12'b000010001011; // 139
storage[4186] =  12'b000001000111; // 71
storage[4187] = -12'b000000100010; // -34
storage[4188] = -12'b000010000001; // -129
storage[4189] =  12'b000010001011; // 139
storage[4190] =  12'b000000010101; // 21
storage[4191] =  12'b000010111010; // 186
storage[4192] =  12'b000000111010; // 58
storage[4193] = -12'b000001101100; // -108
storage[4194] =  12'b000001010011; // 83
storage[4195] = -12'b000000011001; // -25
storage[4196] =  12'b000000000000; // 0
storage[4197] =  12'b000000010101; // 21
storage[4198] = -12'b000001110100; // -116
storage[4199] = -12'b000100000001; // -257
storage[4200] =  12'b000001000011; // 67
storage[4201] =  12'b000001011011; // 91
storage[4202] = -12'b000000001000; // -8
storage[4203] = -12'b000010111001; // -185
storage[4204] = -12'b000001110100; // -116
storage[4205] = -12'b000010100110; // -166
storage[4206] = -12'b000010001111; // -143
storage[4207] =  12'b000000000011; // 3
storage[4208] =  12'b000001010010; // 82
storage[4209] =  12'b000011001011; // 203
storage[4210] = -12'b000001010100; // -84
storage[4211] =  12'b000001000001; // 65
storage[4212] =  12'b000010001101; // 141
storage[4213] =  12'b000000100100; // 36
storage[4214] =  12'b000001010101; // 85
storage[4215] =  12'b000001111000; // 120
storage[4216] = -12'b000100000100; // -260
storage[4217] = -12'b000000100100; // -36
storage[4218] =  12'b000011111011; // 251
storage[4219] = -12'b000010100111; // -167
storage[4220] = -12'b000101010100; // -340
storage[4221] = -12'b000100010110; // -278
storage[4222] = -12'b000011011101; // -221
storage[4223] = -12'b000101010011; // -339
storage[4224] = -12'b000100110011; // -307
storage[4225] = -12'b000001010110; // -86
storage[4226] =  12'b000010001101; // 141
storage[4227] =  12'b000000100001; // 33
storage[4228] =  12'b000000011100; // 28
storage[4229] =  12'b000001001011; // 75
storage[4230] =  12'b000010011101; // 157
storage[4231] =  12'b000000110011; // 51
storage[4232] =  12'b000001100010; // 98
storage[4233] =  12'b000100100000; // 288
storage[4234] = -12'b000010100001; // -161
storage[4235] = -12'b000011101011; // -235
storage[4236] = -12'b000000000111; // -7
storage[4237] =  12'b000100101111; // 303
storage[4238] =  12'b000010100010; // 162
storage[4239] = -12'b000011111100; // -252
storage[4240] =  12'b000001011100; // 92
storage[4241] =  12'b000000001010; // 10
storage[4242] = -12'b000001001010; // -74
storage[4243] = -12'b000000001011; // -11
storage[4244] =  12'b000000101101; // 45
storage[4245] =  12'b000001100011; // 99
storage[4246] = -12'b000100000101; // -261
storage[4247] = -12'b000001100111; // -103
storage[4248] =  12'b000011011011; // 219
storage[4249] =  12'b000000101101; // 45
storage[4250] = -12'b000001001111; // -79
storage[4251] = -12'b000111001110; // -462
storage[4252] = -12'b000101011100; // -348
storage[4253] = -12'b000000010011; // -19
storage[4254] = -12'b000101101000; // -360
storage[4255] = -12'b000001000010; // -66
storage[4256] =  12'b000010111100; // 188
storage[4257] =  12'b000000000101; // 5
storage[4258] =  12'b000000101111; // 47
storage[4259] = -12'b000110110011; // -435
storage[4260] = -12'b001001101110; // -622
storage[4261] =  12'b000010000100; // 132
storage[4262] =  12'b000001011101; // 93
storage[4263] = -12'b000010000101; // -133
storage[4264] =  12'b000000101001; // 41
storage[4265] = -12'b000000010111; // -23
storage[4266] =  12'b000000011101; // 29
storage[4267] =  12'b000001000111; // 71
storage[4268] =  12'b000010110100; // 180
storage[4269] =  12'b000010111001; // 185
storage[4270] =  12'b000010000001; // 129
storage[4271] =  12'b000010101010; // 170
storage[4272] =  12'b000010111011; // 187
storage[4273] =  12'b000000101111; // 47
storage[4274] = -12'b000001011000; // -88
storage[4275] = -12'b000001110110; // -118
storage[4276] = -12'b000010011010; // -154
storage[4277] = -12'b000101001000; // -328
storage[4278] = -12'b000011000001; // -193
storage[4279] = -12'b000010000010; // -130
storage[4280] = -12'b000100001001; // -265
storage[4281] =  12'b000000010010; // 18
storage[4282] =  12'b000000111110; // 62
storage[4283] = -12'b000100100000; // -288
storage[4284] =  12'b000011001111; // 207
storage[4285] = -12'b000001000111; // -71
storage[4286] = -12'b000001011111; // -95
storage[4287] = -12'b000000000010; // -2
storage[4288] = -12'b000000101010; // -42
storage[4289] =  12'b000000111010; // 58
storage[4290] =  12'b000000010111; // 23
storage[4291] =  12'b000000110111; // 55
storage[4292] =  12'b000100000011; // 259
storage[4293] = -12'b000000111010; // -58
storage[4294] =  12'b000001100110; // 102
storage[4295] =  12'b000000011011; // 27
storage[4296] = -12'b000000101000; // -40
storage[4297] = -12'b000010001110; // -142
storage[4298] = -12'b000000111001; // -57
storage[4299] =  12'b000010000001; // 129
storage[4300] = -12'b000010011111; // -159
storage[4301] = -12'b000011000100; // -196
storage[4302] = -12'b001100000000; // -768
storage[4303] =  12'b000110011001; // 409
storage[4304] =  12'b000100010001; // 273
storage[4305] =  12'b000011100000; // 224
storage[4306] =  12'b000011101111; // 239
storage[4307] =  12'b000001010001; // 81
storage[4308] =  12'b000110001010; // 394
storage[4309] =  12'b000000101000; // 40
storage[4310] =  12'b000000101100; // 44
storage[4311] =  12'b000010001100; // 140
storage[4312] =  12'b000010110001; // 177
storage[4313] = -12'b000001100001; // -97
storage[4314] = -12'b000011010000; // -208
storage[4315] =  12'b000000011011; // 27
storage[4316] =  12'b000001000001; // 65
storage[4317] =  12'b000001110100; // 116
storage[4318] = -12'b000000100110; // -38
storage[4319] =  12'b000010001101; // 141
storage[4320] = -12'b000010000111; // -135
storage[4321] = -12'b000000011100; // -28
storage[4322] =  12'b000001000011; // 67
storage[4323] =  12'b000011000110; // 198
storage[4324] = -12'b000000001001; // -9
storage[4325] =  12'b000001100010; // 98
storage[4326] =  12'b000000110010; // 50
storage[4327] = -12'b000001001000; // -72
storage[4328] =  12'b000000011011; // 27
storage[4329] =  12'b000101000111; // 327
storage[4330] =  12'b000010010100; // 148
storage[4331] =  12'b000001100010; // 98
storage[4332] = -12'b000001111101; // -125
storage[4333] = -12'b000001000010; // -66
storage[4334] =  12'b000000100001; // 33
storage[4335] = -12'b000000110001; // -49
storage[4336] =  12'b000001001000; // 72
storage[4337] =  12'b000000101111; // 47
storage[4338] =  12'b000000100101; // 37
storage[4339] = -12'b000010111111; // -191
storage[4340] = -12'b000001101010; // -106
storage[4341] = -12'b000011110000; // -240
storage[4342] =  12'b000011011010; // 218
storage[4343] =  12'b000100110011; // 307
storage[4344] = -12'b000000111111; // -63
storage[4345] =  12'b000001001010; // 74
storage[4346] =  12'b000001010001; // 81
storage[4347] = -12'b000000111001; // -57
storage[4348] =  12'b000010010001; // 145
storage[4349] = -12'b000001111110; // -126
storage[4350] = -12'b000001010010; // -82
storage[4351] =  12'b000000100101; // 37
storage[4352] =  12'b000010100101; // 165
storage[4353] =  12'b000001000011; // 67
storage[4354] = -12'b000010010100; // -148
storage[4355] =  12'b000010000111; // 135
storage[4356] =  12'b000100100001; // 289
storage[4357] =  12'b000010001100; // 140
storage[4358] = -12'b000000000111; // -7
storage[4359] =  12'b000001011010; // 90
storage[4360] = -12'b000000010001; // -17
storage[4361] =  12'b000010100110; // 166
storage[4362] = -12'b000001001110; // -78
storage[4363] = -12'b000001101001; // -105
storage[4364] = -12'b000001001011; // -75
storage[4365] =  12'b000000111010; // 58
storage[4366] =  12'b000011010001; // 209
storage[4367] =  12'b000011010010; // 210
storage[4368] =  12'b000000000101; // 5
storage[4369] = -12'b000001010010; // -82
storage[4370] = -12'b000001100011; // -99
storage[4371] = -12'b000100110010; // -306
storage[4372] = -12'b000010010100; // -148
storage[4373] = -12'b000011100011; // -227
storage[4374] = -12'b000001000101; // -69
storage[4375] =  12'b000010001000; // 136
storage[4376] =  12'b000000101111; // 47
storage[4377] =  12'b000000100110; // 38
storage[4378] = -12'b000011001001; // -201
storage[4379] = -12'b000001100010; // -98
storage[4380] =  12'b000010101100; // 172
storage[4381] = -12'b000011001000; // -200
storage[4382] = -12'b000011001010; // -202
storage[4383] =  12'b000001000101; // 69
storage[4384] =  12'b000010001001; // 137
storage[4385] =  12'b000001010001; // 81
storage[4386] =  12'b000010100001; // 161
storage[4387] =  12'b000000001100; // 12
storage[4388] = -12'b000001011010; // -90
storage[4389] = -12'b000010001010; // -138
storage[4390] = -12'b000001100011; // -99
storage[4391] = -12'b000000010110; // -22
storage[4392] = -12'b000010100110; // -166
storage[4393] =  12'b000001010101; // 85
storage[4394] =  12'b000000001011; // 11
storage[4395] = -12'b000010100011; // -163
storage[4396] = -12'b000010101010; // -170
storage[4397] = -12'b000011000011; // -195
storage[4398] =  12'b000001110100; // 116
storage[4399] = -12'b000001010100; // -84
storage[4400] =  12'b000000100101; // 37
storage[4401] =  12'b000000000111; // 7
storage[4402] = -12'b000000110010; // -50
storage[4403] =  12'b000000100010; // 34
storage[4404] =  12'b000010000111; // 135
storage[4405] =  12'b000001001000; // 72
storage[4406] = -12'b000001010000; // -80
storage[4407] =  12'b000000111001; // 57
storage[4408] =  12'b000000001100; // 12
storage[4409] = -12'b000100110110; // -310
storage[4410] = -12'b000110011111; // -415
storage[4411] =  12'b000000110011; // 51
storage[4412] =  12'b000001011110; // 94
storage[4413] =  12'b000001000100; // 68
storage[4414] =  12'b000001010110; // 86
storage[4415] =  12'b000001001100; // 76
storage[4416] =  12'b000011000000; // 192
storage[4417] =  12'b000010011001; // 153
storage[4418] =  12'b000011100100; // 228
storage[4419] =  12'b000011111010; // 250
storage[4420] = -12'b000110100001; // -417
storage[4421] = -12'b000001100101; // -101
storage[4422] =  12'b000001011011; // 91
storage[4423] = -12'b000010111100; // -188
storage[4424] = -12'b000100110010; // -306
storage[4425] = -12'b000010011110; // -158
storage[4426] = -12'b000011110110; // -246
storage[4427] = -12'b000110001000; // -392
storage[4428] = -12'b000100101010; // -298
storage[4429] = -12'b000000001001; // -9
storage[4430] = -12'b000001101111; // -111
storage[4431] = -12'b000010110001; // -177
storage[4432] = -12'b000001011110; // -94
storage[4433] = -12'b000010011000; // -152
storage[4434] = -12'b000001101010; // -106
storage[4435] =  12'b000000001011; // 11
storage[4436] =  12'b000000110101; // 53
storage[4437] =  12'b000001000000; // 64
storage[4438] = -12'b000001101001; // -105
storage[4439] = -12'b000011100010; // -226
storage[4440] =  12'b000000100011; // 35
storage[4441] = -12'b000010011011; // -155
storage[4442] = -12'b000010101000; // -168
storage[4443] = -12'b000010101000; // -168
storage[4444] = -12'b000000110101; // -53
storage[4445] =  12'b000001000100; // 68
storage[4446] = -12'b000001001000; // -72
storage[4447] =  12'b001000100010; // 546
storage[4448] =  12'b000101010101; // 341
storage[4449] =  12'b000001110011; // 115
storage[4450] =  12'b000100110101; // 309
storage[4451] =  12'b000010010111; // 151
storage[4452] =  12'b000000111010; // 58
storage[4453] =  12'b000010010011; // 147
storage[4454] = -12'b000001110000; // -112
storage[4455] = -12'b000100111000; // -312
storage[4456] = -12'b000010001000; // -136
storage[4457] = -12'b000000101111; // -47
storage[4458] = -12'b000000010110; // -22
storage[4459] =  12'b000001011001; // 89
storage[4460] =  12'b000000110001; // 49
storage[4461] =  12'b000000101011; // 43
storage[4462] =  12'b000000001110; // 14
storage[4463] = -12'b000000010100; // -20
storage[4464] =  12'b000010001110; // 142
storage[4465] = -12'b000100010000; // -272
storage[4466] =  12'b000001010001; // 81
storage[4467] =  12'b000100110110; // 310
storage[4468] = -12'b000011011001; // -217
storage[4469] =  12'b000001111010; // 122
storage[4470] =  12'b000001101111; // 111
storage[4471] = -12'b000011110101; // -245
storage[4472] =  12'b000000101000; // 40
storage[4473] =  12'b000001010101; // 85
storage[4474] = -12'b000001010010; // -82
storage[4475] =  12'b000000000110; // 6
storage[4476] = -12'b000010100000; // -160
storage[4477] =  12'b000000110001; // 49
storage[4478] =  12'b000010111101; // 189
storage[4479] =  12'b000000111111; // 63
storage[4480] =  12'b000000101110; // 46
storage[4481] = -12'b000001011000; // -88
storage[4482] =  12'b000010001000; // 136
storage[4483] = -12'b000011011010; // -218
storage[4484] = -12'b000001111110; // -126
storage[4485] = -12'b000011000101; // -197
storage[4486] =  12'b000010101111; // 175
storage[4487] = -12'b000000100100; // -36
storage[4488] = -12'b000001101111; // -111
storage[4489] =  12'b000101001010; // 330
storage[4490] =  12'b000001110000; // 112
storage[4491] =  12'b000000111101; // 61
storage[4492] =  12'b000010011110; // 158
storage[4493] =  12'b000000001110; // 14
storage[4494] = -12'b000100110100; // -308
storage[4495] =  12'b000000101100; // 44
storage[4496] = -12'b000010001101; // -141
storage[4497] =  12'b000000010000; // 16
storage[4498] = -12'b000000011110; // -30
storage[4499] = -12'b000001000001; // -65
storage[4500] =  12'b000000110011; // 51
storage[4501] =  12'b000000011111; // 31
storage[4502] = -12'b000001100111; // -103
storage[4503] = -12'b000011001000; // -200
storage[4504] =  12'b000000010000; // 16
storage[4505] = -12'b000000000001; // -1
storage[4506] = -12'b000001000111; // -71
storage[4507] =  12'b000001101000; // 104
storage[4508] = -12'b000001010101; // -85
storage[4509] = -12'b000001001101; // -77
storage[4510] =  12'b000001011000; // 88
storage[4511] = -12'b000001111101; // -125
storage[4512] = -12'b000011010100; // -212
storage[4513] = -12'b000000001111; // -15
storage[4514] =  12'b000001111011; // 123
storage[4515] =  12'b000011011001; // 217
storage[4516] =  12'b000000101011; // 43
storage[4517] = -12'b000000101011; // -43
storage[4518] =  12'b000011010110; // 214
storage[4519] =  12'b000000100111; // 39
storage[4520] =  12'b000010011101; // 157
storage[4521] =  12'b000011110100; // 244
storage[4522] =  12'b000000010111; // 23
storage[4523] =  12'b000000010101; // 21
storage[4524] =  12'b000000111001; // 57
storage[4525] = -12'b000100001010; // -266
storage[4526] = -12'b000100001000; // -264
storage[4527] = -12'b000000101000; // -40
storage[4528] = -12'b000101110101; // -373
storage[4529] =  12'b000000110101; // 53
storage[4530] =  12'b000100001000; // 264
storage[4531] = -12'b000010000110; // -134
storage[4532] =  12'b000000111111; // 63
storage[4533] =  12'b000010000010; // 130
storage[4534] =  12'b000010110001; // 177
storage[4535] = -12'b000000010101; // -21
storage[4536] = -12'b000010001000; // -136
storage[4537] =  12'b000001101010; // 106
storage[4538] = -12'b000101001110; // -334
storage[4539] = -12'b000101000100; // -324
storage[4540] =  12'b000001101111; // 111
storage[4541] = -12'b000011101111; // -239
storage[4542] =  12'b000001011010; // 90
storage[4543] =  12'b000000010101; // 21
storage[4544] = -12'b000000101111; // -47
storage[4545] =  12'b000011011011; // 219
storage[4546] = -12'b000010011100; // -156
storage[4547] = -12'b000011001000; // -200
storage[4548] = -12'b000001000010; // -66
storage[4549] =  12'b000000011010; // 26
storage[4550] =  12'b000000110010; // 50
storage[4551] = -12'b000000001011; // -11
storage[4552] =  12'b000101000110; // 326
storage[4553] = -12'b000000010111; // -23
storage[4554] = -12'b000001011100; // -92
storage[4555] =  12'b000010100110; // 166
storage[4556] =  12'b000011111100; // 252
storage[4557] = -12'b000000010011; // -19
storage[4558] = -12'b000001100001; // -97
storage[4559] =  12'b000000100100; // 36
storage[4560] =  12'b000000000101; // 5
storage[4561] = -12'b000100101110; // -302
storage[4562] = -12'b000010011000; // -152
storage[4563] = -12'b000000001011; // -11
storage[4564] = -12'b000000000110; // -6
storage[4565] = -12'b000010111111; // -191
storage[4566] =  12'b000011010001; // 209
storage[4567] =  12'b000000000111; // 7
storage[4568] =  12'b000000100001; // 33
storage[4569] =  12'b000001111011; // 123
storage[4570] = -12'b000001010001; // -81
storage[4571] = -12'b000111000100; // -452
storage[4572] = -12'b000010100100; // -164
storage[4573] =  12'b000010000000; // 128
storage[4574] =  12'b000010111101; // 189
storage[4575] =  12'b000011011000; // 216
storage[4576] = -12'b000011001000; // -200
storage[4577] =  12'b000001011111; // 95
storage[4578] =  12'b000010010001; // 145
storage[4579] = -12'b000010111110; // -190
storage[4580] = -12'b000010011000; // -152
storage[4581] = -12'b000100111011; // -315
storage[4582] = -12'b000000011100; // -28
storage[4583] = -12'b000001011100; // -92
storage[4584] = -12'b000010111101; // -189
storage[4585] = -12'b000100011010; // -282
storage[4586] = -12'b000010010101; // -149
storage[4587] = -12'b000100001101; // -269
storage[4588] = -12'b000010100001; // -161
storage[4589] = -12'b000010011000; // -152
storage[4590] =  12'b000001011100; // 92
storage[4591] = -12'b000010110101; // -181
storage[4592] = -12'b000000111001; // -57
storage[4593] =  12'b000001110001; // 113
storage[4594] = -12'b000000010000; // -16
storage[4595] =  12'b000001001101; // 77
storage[4596] = -12'b000001100110; // -102
storage[4597] = -12'b000001001100; // -76
storage[4598] =  12'b000010010111; // 151
storage[4599] = -12'b000000011100; // -28
storage[4600] =  12'b000001001101; // 77
storage[4601] = -12'b000001001111; // -79
storage[4602] = -12'b000001110010; // -114
storage[4603] =  12'b000001000101; // 69
storage[4604] = -12'b000001100110; // -102
storage[4605] = -12'b000010110011; // -179
storage[4606] =  12'b000010001001; // 137
storage[4607] =  12'b000001100010; // 98
storage[4608] =  12'b000001000110; // 70
storage[4609] = -12'b000001010011; // -83
storage[4610] =  12'b000100111100; // 316
storage[4611] =  12'b000010001110; // 142
storage[4612] = -12'b000001010000; // -80
storage[4613] =  12'b000010111001; // 185
storage[4614] = -12'b000001111000; // -120
storage[4615] =  12'b000010101101; // 173
storage[4616] =  12'b000100000110; // 262
storage[4617] = -12'b000000110011; // -51
storage[4618] =  12'b000010100101; // 165
storage[4619] = -12'b000000010011; // -19
storage[4620] = -12'b000000110101; // -53
storage[4621] =  12'b000000001100; // 12
storage[4622] = -12'b000010101100; // -172
storage[4623] =  12'b000000001111; // 15
storage[4624] = -12'b000100001100; // -268
storage[4625] =  12'b000000100001; // 33
storage[4626] = -12'b000011111111; // -255
storage[4627] = -12'b000000101110; // -46
storage[4628] = -12'b000000001100; // -12
storage[4629] = -12'b000001101100; // -108
storage[4630] =  12'b000001000000; // 64
storage[4631] =  12'b000010011101; // 157
storage[4632] = -12'b000000101000; // -40
storage[4633] =  12'b000001011000; // 88
storage[4634] =  12'b000000111010; // 58
storage[4635] = -12'b000101000100; // -324
storage[4636] = -12'b000010010111; // -151
storage[4637] =  12'b000010010100; // 148
storage[4638] =  12'b000001010001; // 81
storage[4639] = -12'b000010100111; // -167
storage[4640] = -12'b000000100111; // -39
storage[4641] = -12'b000010000001; // -129
storage[4642] = -12'b000100111101; // -317
storage[4643] = -12'b000010001110; // -142
storage[4644] = -12'b000000110101; // -53
storage[4645] =  12'b000010111100; // 188
storage[4646] =  12'b000001110010; // 114
storage[4647] =  12'b000001011111; // 95
storage[4648] =  12'b000011011100; // 220
storage[4649] =  12'b000010010100; // 148
storage[4650] =  12'b000100011110; // 286
storage[4651] = -12'b000000000101; // -5
storage[4652] =  12'b000001011001; // 89
storage[4653] =  12'b000000101110; // 46
storage[4654] =  12'b000011000000; // 192
storage[4655] = -12'b000001010000; // -80
storage[4656] =  12'b000010001011; // 139
storage[4657] =  12'b000001011100; // 92
storage[4658] =  12'b000001011001; // 89
storage[4659] =  12'b000100001101; // 269
storage[4660] =  12'b000000000000; // 0
storage[4661] = -12'b000001000011; // -67
storage[4662] =  12'b000011100010; // 226
storage[4663] = -12'b000101110000; // -368
storage[4664] = -12'b001001001010; // -586
storage[4665] = -12'b000011010111; // -215
storage[4666] = -12'b000101110000; // -368
storage[4667] = -12'b000110101010; // -426
storage[4668] =  12'b000000010111; // 23
storage[4669] = -12'b001100011100; // -796
storage[4670] = -12'b000001001000; // -72
storage[4671] =  12'b000011000101; // 197
storage[4672] = -12'b000000001000; // -8
storage[4673] = -12'b000000101100; // -44
storage[4674] = -12'b000001011111; // -95
storage[4675] =  12'b000001000110; // 70
storage[4676] =  12'b000010100111; // 167
storage[4677] =  12'b000100000010; // 258
storage[4678] =  12'b000010010001; // 145
storage[4679] =  12'b000100011001; // 281
storage[4680] = -12'b000000010001; // -17
storage[4681] = -12'b000001000001; // -65
storage[4682] = -12'b000011101101; // -237
storage[4683] =  12'b000010001100; // 140
storage[4684] = -12'b000010001110; // -142
storage[4685] =  12'b000000100011; // 35
storage[4686] =  12'b000100100100; // 292
storage[4687] = -12'b000001000101; // -69
storage[4688] = -12'b000100111011; // -315
storage[4689] = -12'b000100110000; // -304
storage[4690] =  12'b000000000101; // 5
storage[4691] = -12'b000101101100; // -364
storage[4692] =  12'b000000101011; // 43
storage[4693] =  12'b000000101101; // 45
storage[4694] =  12'b000000010011; // 19
storage[4695] =  12'b000010101011; // 171
storage[4696] =  12'b000011100011; // 227
storage[4697] =  12'b000001111101; // 125
storage[4698] =  12'b000001110011; // 115
storage[4699] = -12'b000011101100; // -236
storage[4700] =  12'b000000000010; // 2
storage[4701] =  12'b000001011101; // 93
storage[4702] = -12'b000011001010; // -202
storage[4703] = -12'b000010100000; // -160
storage[4704] =  12'b000000000011; // 3
storage[4705] = -12'b000011011000; // -216
storage[4706] = -12'b000110010001; // -401
storage[4707] = -12'b001011010110; // -726
storage[4708] =  12'b000000101000; // 40
storage[4709] = -12'b000001110101; // -117
storage[4710] = -12'b000001010000; // -80
storage[4711] = -12'b000011001011; // -203
storage[4712] = -12'b000100111010; // -314
storage[4713] = -12'b000001110011; // -115
storage[4714] =  12'b000001110110; // 118
storage[4715] = -12'b000000010001; // -17
storage[4716] =  12'b000001111011; // 123
storage[4717] = -12'b000010001011; // -139
storage[4718] = -12'b000011001100; // -204
storage[4719] = -12'b000000001101; // -13
storage[4720] = -12'b000011001001; // -201
storage[4721] = -12'b000011010010; // -210
storage[4722] =  12'b000000101111; // 47
storage[4723] = -12'b000001011110; // -94
storage[4724] =  12'b000000001111; // 15
storage[4725] = -12'b000010011101; // -157
storage[4726] =  12'b000011011011; // 219
storage[4727] = -12'b000100001100; // -268
storage[4728] = -12'b000101100101; // -357
storage[4729] = -12'b000010111101; // -189
storage[4730] = -12'b000000110001; // -49
storage[4731] =  12'b000100000010; // 258
storage[4732] = -12'b000000110101; // -53
storage[4733] =  12'b000010101101; // 173
storage[4734] =  12'b000011101110; // 238
storage[4735] =  12'b000011100110; // 230
storage[4736] =  12'b000010011111; // 159
storage[4737] = -12'b000000110001; // -49
storage[4738] =  12'b000011101110; // 238
storage[4739] =  12'b000001011100; // 92
storage[4740] = -12'b000001101011; // -107
storage[4741] =  12'b000000011011; // 27
storage[4742] =  12'b000100100000; // 288
storage[4743] =  12'b000001010001; // 81
storage[4744] =  12'b000010001100; // 140
storage[4745] =  12'b000000001100; // 12
storage[4746] =  12'b000010001001; // 137
storage[4747] =  12'b000011001010; // 202
storage[4748] = -12'b000000001001; // -9
storage[4749] = -12'b000000010111; // -23
storage[4750] = -12'b000000111100; // -60
storage[4751] =  12'b000010011101; // 157
storage[4752] = -12'b000000010000; // -16
storage[4753] =  12'b000000010001; // 17
storage[4754] =  12'b000001011000; // 88
storage[4755] = -12'b000000100010; // -34
storage[4756] =  12'b000010001110; // 142
storage[4757] =  12'b000010000110; // 134
storage[4758] = -12'b000001001001; // -73
storage[4759] = -12'b000001011010; // -90
storage[4760] = -12'b000000001000; // -8
storage[4761] = -12'b000101000110; // -326
storage[4762] =  12'b000010000111; // 135
storage[4763] = -12'b000001011000; // -88
storage[4764] =  12'b000000111010; // 58
storage[4765] = -12'b000011000000; // -192
storage[4766] = -12'b000110010000; // -400
storage[4767] = -12'b000110000000; // -384
storage[4768] = -12'b000001100110; // -102
storage[4769] = -12'b001001110000; // -624
storage[4770] = -12'b001110111100; // -956
storage[4771] =  12'b000001000101; // 69
storage[4772] =  12'b000000000100; // 4
storage[4773] =  12'b000001101100; // 108
storage[4774] =  12'b000101101010; // 362
storage[4775] =  12'b000000111001; // 57
storage[4776] = -12'b000011000000; // -192
storage[4777] =  12'b000001100100; // 100
storage[4778] =  12'b000010101100; // 172
storage[4779] =  12'b000000011101; // 29
storage[4780] =  12'b000011010011; // 211
storage[4781] = -12'b000000000001; // -1
storage[4782] =  12'b000000011110; // 30
storage[4783] =  12'b000000110111; // 55
storage[4784] =  12'b000010101001; // 169
storage[4785] =  12'b000010100011; // 163
storage[4786] = -12'b000000110100; // -52
storage[4787] = -12'b000001010101; // -85
storage[4788] = -12'b000001000110; // -70
storage[4789] =  12'b000000111000; // 56
storage[4790] = -12'b000011110110; // -246
storage[4791] = -12'b000010110001; // -177
storage[4792] =  12'b000011100110; // 230
storage[4793] = -12'b000010000000; // -128
storage[4794] = -12'b000000111001; // -57
storage[4795] =  12'b000000000001; // 1
storage[4796] = -12'b000011100110; // -230
storage[4797] = -12'b000010000011; // -131
storage[4798] = -12'b000001010111; // -87
storage[4799] =  12'b000011011110; // 222
storage[4800] =  12'b000101001011; // 331
storage[4801] = -12'b000010110001; // -177
storage[4802] =  12'b000001111101; // 125
storage[4803] = -12'b000000000100; // -4
storage[4804] = -12'b000111010000; // -464
storage[4805] = -12'b000000111010; // -58
storage[4806] = -12'b000001011100; // -92
storage[4807] = -12'b000011001111; // -207
storage[4808] = -12'b000100000111; // -263
storage[4809] = -12'b000011010001; // -209
storage[4810] = -12'b000011101000; // -232
storage[4811] = -12'b000011101000; // -232
storage[4812] =  12'b000000100100; // 36
storage[4813] = -12'b000110001101; // -397
storage[4814] =  12'b000001011101; // 93
storage[4815] =  12'b000000101110; // 46
storage[4816] =  12'b000010000101; // 133
storage[4817] =  12'b000100000001; // 257
storage[4818] =  12'b000100110110; // 310
storage[4819] =  12'b000000001010; // 10
storage[4820] = -12'b000000010101; // -21
storage[4821] =  12'b000010111000; // 184
storage[4822] =  12'b000000010001; // 17
storage[4823] =  12'b000000111110; // 62
storage[4824] = -12'b001000100101; // -549
storage[4825] = -12'b000101000101; // -325
storage[4826] = -12'b000010001101; // -141
storage[4827] =  12'b000000000111; // 7
storage[4828] =  12'b000010001001; // 137
storage[4829] =  12'b000100110111; // 311
storage[4830] = -12'b000000111010; // -58
storage[4831] = -12'b000010110000; // -176
storage[4832] = -12'b000011101011; // -235
storage[4833] = -12'b000010111110; // -190
storage[4834] = -12'b000010001101; // -141
storage[4835] = -12'b000001110100; // -116
storage[4836] =  12'b000011010011; // 211
storage[4837] =  12'b000010101100; // 172
storage[4838] = -12'b000001010001; // -81
storage[4839] =  12'b000001000101; // 69
storage[4840] =  12'b000000110011; // 51
storage[4841] =  12'b000001101011; // 107
storage[4842] =  12'b000010001110; // 142
storage[4843] = -12'b000000001101; // -13
storage[4844] = -12'b000000010000; // -16
storage[4845] = -12'b000011111111; // -255
storage[4846] = -12'b000001001101; // -77
storage[4847] = -12'b000001111011; // -123
storage[4848] = -12'b000000010110; // -22
storage[4849] = -12'b000000101101; // -45
storage[4850] = -12'b000111010101; // -469
storage[4851] = -12'b000011111011; // -251
storage[4852] = -12'b000000001000; // -8
storage[4853] = -12'b000001100001; // -97
storage[4854] = -12'b000010000001; // -129
storage[4855] = -12'b000000000110; // -6
storage[4856] =  12'b000000111010; // 58
storage[4857] = -12'b000000010001; // -17
storage[4858] = -12'b000001100100; // -100
storage[4859] = -12'b000010100000; // -160
storage[4860] = -12'b000001101111; // -111
storage[4861] =  12'b000001001110; // 78
storage[4862] = -12'b000001110000; // -112
storage[4863] = -12'b000000001001; // -9
storage[4864] = -12'b000000010110; // -22
storage[4865] = -12'b000000110001; // -49
storage[4866] =  12'b000000010110; // 22
storage[4867] = -12'b000001101001; // -105
storage[4868] = -12'b000001010010; // -82
storage[4869] = -12'b000000101110; // -46
storage[4870] = -12'b000001011000; // -88
storage[4871] = -12'b000010100000; // -160
storage[4872] = -12'b000000001100; // -12
storage[4873] = -12'b000000110010; // -50
storage[4874] =  12'b000001011000; // 88
storage[4875] = -12'b000010100101; // -165
storage[4876] =  12'b000000001110; // 14
storage[4877] = -12'b000001111011; // -123
storage[4878] = -12'b000010010100; // -148
storage[4879] = -12'b000000110001; // -49
storage[4880] = -12'b000010000011; // -131
storage[4881] = -12'b000001000110; // -70
storage[4882] = -12'b000000000010; // -2
storage[4883] = -12'b000001110011; // -115
storage[4884] = -12'b000000011011; // -27
storage[4885] = -12'b000000010100; // -20
storage[4886] = -12'b000010000000; // -128
storage[4887] =  12'b000000110011; // 51
storage[4888] =  12'b000000011111; // 31
storage[4889] = -12'b000010011101; // -157
storage[4890] = -12'b000000111101; // -61
storage[4891] = -12'b000010000101; // -133
storage[4892] = -12'b000011000110; // -198
storage[4893] = -12'b000000000100; // -4
storage[4894] = -12'b000000001011; // -11
storage[4895] = -12'b000000011011; // -27
storage[4896] = -12'b000001101100; // -108
storage[4897] = -12'b000010110111; // -183
storage[4898] =  12'b000000100000; // 32
storage[4899] = -12'b000010110010; // -178
storage[4900] =  12'b000001001110; // 78
storage[4901] = -12'b000000011100; // -28
storage[4902] = -12'b000010101100; // -172
storage[4903] = -12'b000000001101; // -13
storage[4904] = -12'b000001100101; // -101
storage[4905] =  12'b000000010010; // 18
storage[4906] =  12'b000000110110; // 54
storage[4907] =  12'b000001001011; // 75
storage[4908] = -12'b000001011011; // -91
storage[4909] =  12'b000001100000; // 96
storage[4910] = -12'b000000000111; // -7
storage[4911] =  12'b000000010001; // 17
storage[4912] = -12'b000010101000; // -168
storage[4913] = -12'b000001000100; // -68
storage[4914] =  12'b000001000100; // 68
storage[4915] =  12'b000000010110; // 22
storage[4916] =  12'b000001001011; // 75
storage[4917] =  12'b000000100110; // 38
storage[4918] = -12'b000001110011; // -115
storage[4919] =  12'b000010000000; // 128
storage[4920] =  12'b000000101011; // 43
storage[4921] =  12'b000001011010; // 90
storage[4922] = -12'b000001111111; // -127
storage[4923] = -12'b000001101010; // -106
storage[4924] = -12'b000001000100; // -68
storage[4925] =  12'b000000000101; // 5
storage[4926] =  12'b000000011010; // 26
storage[4927] = -12'b000001010010; // -82
storage[4928] = -12'b000010001010; // -138
storage[4929] = -12'b000001110000; // -112
storage[4930] = -12'b000010110101; // -181
storage[4931] =  12'b000000010100; // 20
storage[4932] = -12'b000001100001; // -97
storage[4933] = -12'b000000110010; // -50
storage[4934] = -12'b000010111001; // -185
storage[4935] = -12'b000010001111; // -143
storage[4936] =  12'b000000100100; // 36
storage[4937] = -12'b000001110011; // -115
storage[4938] =  12'b000000101101; // 45
storage[4939] = -12'b000000101100; // -44
storage[4940] =  12'b000000100110; // 38
storage[4941] = -12'b000001100010; // -98
storage[4942] =  12'b000000010010; // 18
storage[4943] =  12'b000001001010; // 74
storage[4944] = -12'b000000110001; // -49
storage[4945] = -12'b000010001101; // -141
storage[4946] = -12'b000000000110; // -6
storage[4947] =  12'b000000000110; // 6
storage[4948] =  12'b000000101100; // 44
storage[4949] = -12'b000000011111; // -31
storage[4950] = -12'b000010100011; // -163
storage[4951] =  12'b000000111101; // 61
storage[4952] =  12'b000000100010; // 34
storage[4953] = -12'b000001010010; // -82
storage[4954] = -12'b000001010000; // -80
storage[4955] =  12'b000001001011; // 75
storage[4956] = -12'b000010001010; // -138
storage[4957] = -12'b000000100111; // -39
storage[4958] = -12'b000001010101; // -85
storage[4959] = -12'b000000001111; // -15
storage[4960] = -12'b000010001111; // -143
storage[4961] = -12'b000000001110; // -14
storage[4962] =  12'b000001000100; // 68
storage[4963] = -12'b000010000010; // -130
storage[4964] = -12'b000000111011; // -59
storage[4965] = -12'b000000000011; // -3
storage[4966] =  12'b000001001011; // 75
storage[4967] = -12'b000000111110; // -62
storage[4968] = -12'b000001101100; // -108
storage[4969] = -12'b000001010000; // -80
storage[4970] = -12'b000001000111; // -71
storage[4971] = -12'b000000011010; // -26
storage[4972] = -12'b000001001100; // -76
storage[4973] =  12'b000001011001; // 89
storage[4974] = -12'b000001110000; // -112
storage[4975] = -12'b000001111010; // -122
storage[4976] =  12'b000000111011; // 59
storage[4977] = -12'b000000010011; // -19
storage[4978] = -12'b000001101101; // -109
storage[4979] =  12'b000001000110; // 70
storage[4980] = -12'b000000000111; // -7
storage[4981] =  12'b000001001100; // 76
storage[4982] = -12'b000001110100; // -116
storage[4983] = -12'b000001111100; // -124
storage[4984] = -12'b000001110001; // -113
storage[4985] = -12'b000001110101; // -117
storage[4986] =  12'b000000100001; // 33
storage[4987] = -12'b000000000100; // -4
storage[4988] = -12'b000000111101; // -61
storage[4989] = -12'b000001110110; // -118
storage[4990] = -12'b000001100101; // -101
storage[4991] =  12'b000000001111; // 15
storage[4992] =  12'b000000010100; // 20
storage[4993] = -12'b000010000110; // -134
storage[4994] = -12'b000010001000; // -136
storage[4995] = -12'b000000110010; // -50
storage[4996] = -12'b000011001000; // -200
storage[4997] =  12'b000100001011; // 267
storage[4998] =  12'b000011011100; // 220
storage[4999] = -12'b000011010111; // -215
storage[5000] =  12'b000001000111; // 71
storage[5001] =  12'b000000110100; // 52
storage[5002] =  12'b000001010111; // 87
storage[5003] =  12'b000001001111; // 79
storage[5004] =  12'b000000001010; // 10
storage[5005] = -12'b000010100111; // -167
storage[5006] = -12'b000100001001; // -265
storage[5007] =  12'b000000111111; // 63
storage[5008] = -12'b000011111101; // -253
storage[5009] = -12'b001100110100; // -820
storage[5010] = -12'b000100011000; // -280
storage[5011] = -12'b000100001001; // -265
storage[5012] = -12'b000010001100; // -140
storage[5013] = -12'b000110010100; // -404
storage[5014] = -12'b000010110101; // -181
storage[5015] = -12'b000100001001; // -265
storage[5016] = -12'b000010000010; // -130
storage[5017] =  12'b000000000001; // 1
storage[5018] =  12'b000000111011; // 59
storage[5019] =  12'b000000010001; // 17
storage[5020] =  12'b000011001111; // 207
storage[5021] =  12'b000000101101; // 45
storage[5022] = -12'b000010110000; // -176
storage[5023] = -12'b000010000101; // -133
storage[5024] =  12'b000000101000; // 40
storage[5025] =  12'b000010111001; // 185
storage[5026] = -12'b000000011000; // -24
storage[5027] = -12'b000011101111; // -239
storage[5028] = -12'b000000011011; // -27
storage[5029] = -12'b000000110111; // -55
storage[5030] =  12'b000000111000; // 56
storage[5031] = -12'b000010001110; // -142
storage[5032] = -12'b000011100100; // -228
storage[5033] = -12'b000010000011; // -131
storage[5034] =  12'b000100100001; // 289
storage[5035] =  12'b000010100000; // 160
storage[5036] = -12'b000000001101; // -13
storage[5037] =  12'b000001101000; // 104
storage[5038] = -12'b000010000010; // -130
storage[5039] =  12'b000011111110; // 254
storage[5040] =  12'b000011101001; // 233
storage[5041] =  12'b000010111000; // 184
storage[5042] =  12'b000101000101; // 325
storage[5043] = -12'b000010100110; // -166
storage[5044] = -12'b000010111110; // -190
storage[5045] =  12'b000001010000; // 80
storage[5046] = -12'b000110100011; // -419
storage[5047] = -12'b000000001100; // -12
storage[5048] = -12'b000101110010; // -370
storage[5049] = -12'b000110011110; // -414
storage[5050] =  12'b000000001100; // 12
storage[5051] = -12'b000000100011; // -35
storage[5052] = -12'b000000010011; // -19
storage[5053] = -12'b000011111011; // -251
storage[5054] = -12'b000000000011; // -3
storage[5055] =  12'b000000110010; // 50
storage[5056] = -12'b000001110001; // -113
storage[5057] =  12'b000010010010; // 146
storage[5058] = -12'b000001001100; // -76
storage[5059] = -12'b000001110000; // -112
storage[5060] =  12'b000000111111; // 63
storage[5061] = -12'b000010011110; // -158
storage[5062] = -12'b000000100001; // -33
storage[5063] =  12'b000000101001; // 41
storage[5064] =  12'b000000000100; // 4
storage[5065] =  12'b000011010011; // 211
storage[5066] = -12'b000010010010; // -146
storage[5067] = -12'b000010001101; // -141
storage[5068] = -12'b000010110100; // -180
storage[5069] = -12'b000010000101; // -133
storage[5070] = -12'b000110010110; // -406
storage[5071] = -12'b000001011000; // -88
storage[5072] =  12'b000010100000; // 160
storage[5073] =  12'b000000100001; // 33
storage[5074] = -12'b000010001101; // -141
storage[5075] = -12'b000100110010; // -306
storage[5076] = -12'b000110010100; // -404
storage[5077] = -12'b000101011101; // -349
storage[5078] = -12'b000000101111; // -47
storage[5079] = -12'b000000000100; // -4
storage[5080] = -12'b000110000110; // -390
storage[5081] = -12'b000101011110; // -350
storage[5082] = -12'b000001111011; // -123
storage[5083] = -12'b000000110010; // -50
storage[5084] =  12'b000011001111; // 207
storage[5085] = -12'b000000100101; // -37
storage[5086] =  12'b000011000111; // 199
storage[5087] =  12'b000010011100; // 156
storage[5088] = -12'b000000110001; // -49
storage[5089] =  12'b000000110010; // 50
storage[5090] =  12'b000010101101; // 173
storage[5091] =  12'b000010101000; // 168
storage[5092] = -12'b000001011100; // -92
storage[5093] = -12'b000000111110; // -62
storage[5094] = -12'b000111001100; // -460
storage[5095] =  12'b000000111111; // 63
storage[5096] = -12'b000000110110; // -54
storage[5097] =  12'b000001011000; // 88
storage[5098] = -12'b000010100111; // -167
storage[5099] =  12'b000001000100; // 68
storage[5100] = -12'b000011110001; // -241
storage[5101] =  12'b000100011111; // 287
storage[5102] = -12'b000000100001; // -33
storage[5103] =  12'b000000100110; // 38
storage[5104] =  12'b000111000101; // 453
storage[5105] =  12'b000011011110; // 222
storage[5106] =  12'b000000101110; // 46
storage[5107] =  12'b000100110101; // 309
storage[5108] = -12'b000000011110; // -30
storage[5109] = -12'b000111001111; // -463
storage[5110] =  12'b000000100011; // 35
storage[5111] =  12'b000000111100; // 60
storage[5112] =  12'b000000110111; // 55
storage[5113] = -12'b000011001011; // -203
storage[5114] =  12'b000000110110; // 54
storage[5115] =  12'b000010010000; // 144
storage[5116] = -12'b000010011100; // -156
storage[5117] =  12'b000001100101; // 101
storage[5118] =  12'b000000000011; // 3
storage[5119] =  12'b000000111100; // 60
storage[5120] =  12'b000100100111; // 295
storage[5121] =  12'b000011000000; // 192
storage[5122] =  12'b000010011000; // 152
storage[5123] =  12'b000000110011; // 51
storage[5124] = -12'b000010111010; // -186
storage[5125] =  12'b000010000110; // 134
storage[5126] =  12'b000010010101; // 149
storage[5127] =  12'b000011010001; // 209
storage[5128] = -12'b000011100010; // -226
storage[5129] =  12'b000001110011; // 115
storage[5130] =  12'b000011101110; // 238
storage[5131] =  12'b000000101001; // 41
storage[5132] = -12'b000010101011; // -171
storage[5133] = -12'b000111100111; // -487
storage[5134] = -12'b000010000000; // -128
storage[5135] = -12'b000010011001; // -153
storage[5136] = -12'b000100011101; // -285
storage[5137] = -12'b000001110010; // -114
storage[5138] = -12'b000000100011; // -35
storage[5139] =  12'b000000100110; // 38
storage[5140] = -12'b000000100000; // -32
storage[5141] = -12'b000011011010; // -218
storage[5142] = -12'b001011000110; // -710
storage[5143] =  12'b000000001010; // 10
storage[5144] = -12'b000001110101; // -117
storage[5145] = -12'b001000010100; // -532
storage[5146] = -12'b000000001110; // -14
storage[5147] = -12'b000111111111; // -511
storage[5148] = -12'b000001010000; // -80
storage[5149] =  12'b000000101101; // 45
storage[5150] = -12'b000000101110; // -46
storage[5151] = -12'b000011111010; // -250
storage[5152] =  12'b000001011101; // 93
storage[5153] = -12'b000010000110; // -134
storage[5154] = -12'b000001110000; // -112
storage[5155] = -12'b000000011111; // -31
storage[5156] = -12'b000000011010; // -26
storage[5157] = -12'b000000010000; // -16
storage[5158] =  12'b000011011110; // 222
storage[5159] =  12'b000110011110; // 414
storage[5160] = -12'b000100011101; // -285
storage[5161] = -12'b000010000100; // -132
storage[5162] =  12'b000010011101; // 157
storage[5163] = -12'b000101101001; // -361
storage[5164] =  12'b000000111011; // 59
storage[5165] = -12'b000001101001; // -105
storage[5166] = -12'b000110111010; // -442
storage[5167] =  12'b001001010110; // 598
storage[5168] =  12'b000011011101; // 221
storage[5169] =  12'b000000110011; // 51
storage[5170] =  12'b000010010011; // 147
storage[5171] =  12'b000011001100; // 204
storage[5172] =  12'b000011010100; // 212
storage[5173] =  12'b000000100010; // 34
storage[5174] =  12'b000001011100; // 92
storage[5175] =  12'b000011101010; // 234
storage[5176] = -12'b000110000100; // -388
storage[5177] = -12'b000100001111; // -271
storage[5178] = -12'b000000111111; // -63
storage[5179] =  12'b000000100000; // 32
storage[5180] =  12'b000001100001; // 97
storage[5181] =  12'b000001110111; // 119
storage[5182] = -12'b000000001010; // -10
storage[5183] =  12'b000001010100; // 84
storage[5184] =  12'b000001101100; // 108
storage[5185] = -12'b000111010101; // -469
storage[5186] = -12'b000000000100; // -4
storage[5187] =  12'b000000100111; // 39
storage[5188] = -12'b000100001110; // -270
storage[5189] =  12'b000000001010; // 10
storage[5190] =  12'b000000010111; // 23
storage[5191] = -12'b000000011111; // -31
storage[5192] =  12'b000100011101; // 285
storage[5193] =  12'b000010101000; // 168
storage[5194] =  12'b000010001001; // 137
storage[5195] =  12'b000010010000; // 144
storage[5196] =  12'b000011100000; // 224
storage[5197] = -12'b000000111000; // -56
storage[5198] = -12'b000001011010; // -90
storage[5199] = -12'b000101100111; // -359
storage[5200] = -12'b000000001011; // -11
storage[5201] =  12'b000001001001; // 73
storage[5202] = -12'b000000000001; // -1
storage[5203] = -12'b000101101010; // -362
storage[5204] = -12'b000010011100; // -156
storage[5205] = -12'b000010101101; // -173
storage[5206] =  12'b000010011111; // 159
storage[5207] =  12'b000101110100; // 372
storage[5208] =  12'b000010111010; // 186
storage[5209] = -12'b000001100111; // -103
storage[5210] = -12'b000000111111; // -63
storage[5211] =  12'b000000111110; // 62
storage[5212] =  12'b000011100000; // 224
storage[5213] =  12'b000011001011; // 203
storage[5214] =  12'b000011100110; // 230
storage[5215] =  12'b000011100110; // 230
storage[5216] =  12'b000011111101; // 253
storage[5217] =  12'b000010000111; // 135
storage[5218] =  12'b000010101000; // 168
storage[5219] =  12'b000011111100; // 252
storage[5220] =  12'b000010100000; // 160
storage[5221] =  12'b000001111101; // 125
storage[5222] = -12'b000000010100; // -20
storage[5223] = -12'b000001110110; // -118
storage[5224] =  12'b000001001011; // 75
storage[5225] =  12'b000011100000; // 224
storage[5226] = -12'b000010011110; // -158
storage[5227] =  12'b000010010110; // 150
storage[5228] =  12'b000010001010; // 138
storage[5229] =  12'b000011000010; // 194
storage[5230] =  12'b000001000000; // 64
storage[5231] =  12'b000010000110; // 134
storage[5232] =  12'b000111011111; // 479
storage[5233] = -12'b000101101011; // -363
storage[5234] = -12'b001110001111; // -911
storage[5235] = -12'b000011111111; // -255
storage[5236] =  12'b000000100111; // 39
storage[5237] = -12'b000111011101; // -477
storage[5238] =  12'b000011010001; // 209
storage[5239] = -12'b000001010101; // -85
storage[5240] =  12'b000001110101; // 117
storage[5241] = -12'b000010000111; // -135
storage[5242] = -12'b000101101011; // -363
storage[5243] = -12'b000011010100; // -212
storage[5244] = -12'b000100100101; // -293
storage[5245] = -12'b000011011101; // -221
storage[5246] =  12'b000100000001; // 257
storage[5247] =  12'b000001110111; // 119
storage[5248] = -12'b000001101110; // -110
storage[5249] =  12'b000001001000; // 72
storage[5250] =  12'b000001101110; // 110
storage[5251] = -12'b000010000111; // -135
storage[5252] =  12'b000011111001; // 249
storage[5253] =  12'b000100001111; // 271
storage[5254] = -12'b000001110110; // -118
storage[5255] =  12'b000000110110; // 54
storage[5256] =  12'b000000001000; // 8
storage[5257] =  12'b000011100110; // 230
storage[5258] = -12'b000001100111; // -103
storage[5259] = -12'b000000011110; // -30
storage[5260] = -12'b000100000000; // -256
storage[5261] = -12'b001000011100; // -540
storage[5262] = -12'b000100010011; // -275
storage[5263] =  12'b000000011110; // 30
storage[5264] = -12'b000010111001; // -185
storage[5265] =  12'b000011011100; // 220
storage[5266] =  12'b000010110011; // 179
storage[5267] =  12'b000010110000; // 176
storage[5268] = -12'b000111100011; // -483
storage[5269] = -12'b000001001111; // -79
storage[5270] = -12'b000000001011; // -11
storage[5271] = -12'b000110001001; // -393
storage[5272] =  12'b000000100101; // 37
storage[5273] = -12'b000010001110; // -142
storage[5274] =  12'b000010010011; // 147
storage[5275] =  12'b000000101100; // 44
storage[5276] = -12'b000011001111; // -207
storage[5277] = -12'b000011101011; // -235
storage[5278] =  12'b000000111101; // 61
storage[5279] = -12'b000000111101; // -61
storage[5280] =  12'b000010010101; // 149
storage[5281] =  12'b000000001011; // 11
storage[5282] =  12'b000001110000; // 112
storage[5283] =  12'b000000111100; // 60
storage[5284] =  12'b000010010011; // 147
storage[5285] =  12'b000111011011; // 475
storage[5286] =  12'b000010101010; // 170
storage[5287] = -12'b000001100101; // -101
storage[5288] = -12'b001011001111; // -719
storage[5289] = -12'b000000100111; // -39
storage[5290] = -12'b000111101010; // -490
storage[5291] =  12'b000111000010; // 450
storage[5292] =  12'b000100111101; // 317
storage[5293] = -12'b000011111111; // -255
storage[5294] = -12'b000001111101; // -125
storage[5295] = -12'b000101100010; // -354
storage[5296] =  12'b001001000000; // 576
storage[5297] =  12'b001000101000; // 552
storage[5298] = -12'b000000110011; // -51
storage[5299] =  12'b000100010010; // 274
storage[5300] =  12'b000101010111; // 343
storage[5301] =  12'b000010010111; // 151
storage[5302] =  12'b000111101010; // 490
storage[5303] =  12'b000100101111; // 303
storage[5304] = -12'b000001001111; // -79
storage[5305] =  12'b000101111101; // 381
storage[5306] =  12'b000001101000; // 104
storage[5307] =  12'b000010100101; // 165
storage[5308] = -12'b000011100111; // -231
storage[5309] =  12'b000001101000; // 104
storage[5310] = -12'b001101011101; // -861
storage[5311] = -12'b000100101100; // -300
storage[5312] = -12'b000011100100; // -228
storage[5313] =  12'b001001000010; // 578
storage[5314] = -12'b000010010000; // -144
storage[5315] = -12'b000111101110; // -494
storage[5316] =  12'b000011101100; // 236
storage[5317] = -12'b000000101001; // -41
storage[5318] = -12'b000100100111; // -295
storage[5319] = -12'b000000000101; // -5
storage[5320] =  12'b000011100110; // 230
storage[5321] = -12'b000010011011; // -155
storage[5322] =  12'b001010001101; // 653
storage[5323] = -12'b000101110110; // -374
storage[5324] =  12'b001011101110; // 750
storage[5325] = -12'b000110001011; // -395
storage[5326] =  12'b000000111110; // 62
storage[5327] = -12'b001100111100; // -828
storage[5328] = -12'b000001001000; // -72
storage[5329] =  12'b000100011010; // 282
storage[5330] = -12'b000010001111; // -143
storage[5331] = -12'b000000010111; // -23
storage[5332] =  12'b000010110001; // 177
storage[5333] = -12'b000101000100; // -324
storage[5334] =  12'b000110010100; // 404
storage[5335] =  12'b000100010000; // 272
storage[5336] =  12'b000001000000; // 64
storage[5337] = -12'b001010000101; // -645
storage[5338] =  12'b000011101110; // 238
storage[5339] = -12'b001011111011; // -763
storage[5340] =  12'b000101101101; // 365
storage[5341] =  12'b001000011111; // 543
storage[5342] = -12'b000001000000; // -64
storage[5343] =  12'b000100100000; // 288
storage[5344] =  12'b000000100010; // 34
storage[5345] = -12'b000000011111; // -31
storage[5346] =  12'b000100110111; // 311
storage[5347] = -12'b000101011000; // -344
storage[5348] = -12'b000011010011; // -211
storage[5349] = -12'b001101000001; // -833
storage[5350] = -12'b000110010011; // -403
storage[5351] = -12'b000010011001; // -153
storage[5352] = -12'b000111001110; // -462
storage[5353] =  12'b000101110101; // 373
storage[5354] =  12'b000011100110; // 230
storage[5355] = -12'b000101001100; // -332
storage[5356] = -12'b000000001011; // -11
storage[5357] =  12'b000100111010; // 314
storage[5358] = -12'b001001010111; // -599
storage[5359] =  12'b000001001111; // 79
storage[5360] = -12'b001011000100; // -708
storage[5361] = -12'b000111010000; // -464
storage[5362] = -12'b000100111110; // -318
storage[5363] =  12'b001100100111; // 807
storage[5364] = -12'b000100100010; // -290
storage[5365] = -12'b000010001100; // -140
storage[5366] = -12'b000010101010; // -170
storage[5367] = -12'b010000010100; // -1044
storage[5368] = -12'b001010010110; // -662
storage[5369] = -12'b000110010001; // -401
storage[5370] = -12'b000001010100; // -84
storage[5371] =  12'b000101110110; // 374
storage[5372] =  12'b001000101000; // 552
storage[5373] =  12'b001011110100; // 756
storage[5374] = -12'b000001100000; // -96
storage[5375] =  12'b000001110001; // 113
storage[5376] =  12'b000000011000; // 24
storage[5377] = -12'b000001000100; // -68
storage[5378] =  12'b001000101011; // 555
storage[5379] = -12'b000000011010; // -26
storage[5380] =  12'b000101111111; // 383
storage[5381] = -12'b000011010001; // -209
storage[5382] = -12'b000000110111; // -55
storage[5383] = -12'b001001010000; // -592
storage[5384] = -12'b001001010110; // -598
storage[5385] = -12'b000101111110; // -382
storage[5386] =  12'b000111010010; // 466
storage[5387] =  12'b000111100001; // 481
storage[5388] = -12'b000101100001; // -353
storage[5389] =  12'b000101111101; // 381
storage[5390] =  12'b000101100111; // 359
storage[5391] = -12'b001010110111; // -695
storage[5392] =  12'b000011000000; // 192
storage[5393] = -12'b000000011100; // -28
storage[5394] =  12'b000101111110; // 382
storage[5395] =  12'b000010110110; // 182
storage[5396] = -12'b001011111100; // -764
storage[5397] = -12'b000011110101; // -245
storage[5398] =  12'b000011111010; // 250
storage[5399] =  12'b000011110100; // 244
storage[5400] =  12'b000011100111; // 231
storage[5401] =  12'b000100000000; // 256
storage[5402] = -12'b000001100001; // -97
storage[5403] = -12'b000001001111; // -79
storage[5404] =  12'b000111001001; // 457
storage[5405] = -12'b000010101101; // -173
storage[5406] =  12'b000100110001; // 305
storage[5407] =  12'b000001110011; // 115
storage[5408] = -12'b001111001010; // -970
storage[5409] =  12'b000100111110; // 318
storage[5410] = -12'b000011011001; // -217
storage[5411] = -12'b000100001111; // -271
storage[5412] = -12'b000011011110; // -222
storage[5413] = -12'b000010111011; // -187
storage[5414] = -12'b000011001010; // -202
storage[5415] = -12'b000101011011; // -347
storage[5416] =  12'b000110010101; // 405
storage[5417] = -12'b000010010110; // -150
storage[5418] = -12'b000001010010; // -82
storage[5419] = -12'b000000111111; // -63
storage[5420] = -12'b000011011101; // -221
storage[5421] =  12'b000111111101; // 509
storage[5422] = -12'b000011000011; // -195
storage[5423] = -12'b001000110101; // -565
storage[5424] =  12'b000000110011; // 51
storage[5425] =  12'b000111011100; // 476
storage[5426] =  12'b000110100100; // 420
storage[5427] =  12'b000010010101; // 149
storage[5428] = -12'b000101111011; // -379
storage[5429] =  12'b000010000001; // 129
storage[5430] = -12'b000100111100; // -316
storage[5431] = -12'b000001000100; // -68
storage[5432] = -12'b000110110001; // -433
storage[5433] =  12'b000010010010; // 146
storage[5434] = -12'b000111000011; // -451
storage[5435] = -12'b000010010000; // -144
storage[5436] =  12'b000000101000; // 40
storage[5437] =  12'b000101111101; // 381
storage[5438] =  12'b000010010011; // 147
storage[5439] =  12'b000011011110; // 222
storage[5440] = -12'b001100001101; // -781
storage[5441] =  12'b000010001010; // 138
storage[5442] =  12'b000001100101; // 101
storage[5443] =  12'b001000011000; // 536
storage[5444] = -12'b001010011011; // -667
storage[5445] = -12'b001000001110; // -526
storage[5446] = -12'b000100110010; // -306
storage[5447] = -12'b010100011111; // -1311
storage[5448] = -12'b000101000000; // -320
storage[5449] =  12'b001110111011; // 955
storage[5450] =  12'b001011000001; // 705
storage[5451] = -12'b011101000110; // -1862
storage[5452] =  12'b000001111010; // 122
storage[5453] = -12'b000001111101; // -125
storage[5454] =  12'b000011100100; // 228
storage[5455] = -12'b010100001101; // -1293
storage[5456] =  12'b000001000110; // 70
storage[5457] = -12'b000101001010; // -330
storage[5458] =  12'b010101001111; // 1359
storage[5459] = -12'b000100011010; // -282
end

always @(posedge clk) if (we==1) storage[address_p] <= dp;
always @(posedge clk) if (re==1) datata<=storage[address];

endmodule
