module database(clk,datata,re,address,we,dp,address_p);

parameter SIZE=13;

input clk;
output reg signed [SIZE-1:0] datata;
input re,we;
input [14:0] address;
input signed [SIZE-1:0] dp;
input [14:0] address_p;

reg signed [SIZE-1:0] storage [5459:0];

initial begin

storage[0] =  12'b100111100000; // [ 0.6171875]
storage[1] =  12'b100111110000; // [ 0.62109375]
storage[2] =  12'b101000000000; // [ 0.625]
storage[3] =  12'b101000100000; // [ 0.6328125]
storage[4] =  12'b101000110000; // [ 0.63671875]
storage[5] =  12'b101000110000; // [ 0.63671875]
storage[6] =  12'b101000010000; // [ 0.62890625]
storage[7] =  12'b100110100000; // [ 0.6015625]
storage[8] =  12'b100010110000; // [ 0.54296875]
storage[9] =  12'b011110110000; // [ 0.48046875]
storage[10] =  12'b011010110000; // [ 0.41796875]
storage[11] =  12'b011001000000; // [ 0.390625]
storage[12] =  12'b011000110000; // [ 0.38671875]
storage[13] =  12'b011010000000; // [ 0.40625]
storage[14] =  12'b011100000000; // [ 0.4375]
storage[15] =  12'b100000010000; // [ 0.50390625]
storage[16] =  12'b100101010000; // [ 0.58203125]
storage[17] =  12'b101000010000; // [ 0.62890625]
storage[18] =  12'b101001010000; // [ 0.64453125]
storage[19] =  12'b101001010000; // [ 0.64453125]
storage[20] =  12'b101001100000; // [ 0.6484375]
storage[21] =  12'b101001000000; // [ 0.640625]
storage[22] =  12'b101001000000; // [ 0.640625]
storage[23] =  12'b101000110000; // [ 0.63671875]
storage[24] =  12'b101000100000; // [ 0.6328125]
storage[25] =  12'b101000010000; // [ 0.62890625]
storage[26] =  12'b101000000000; // [ 0.625]
storage[27] =  12'b100111100000; // [ 0.6171875]
storage[28] =  12'b100111010000; // [ 0.61328125]
storage[29] =  12'b100111110000; // [ 0.62109375]
storage[30] =  12'b101000000000; // [ 0.625]
storage[31] =  12'b101000100000; // [ 0.6328125]
storage[32] =  12'b101000110000; // [ 0.63671875]
storage[33] =  12'b101000010000; // [ 0.62890625]
storage[34] =  12'b100101100000; // [ 0.5859375]
storage[35] =  12'b011100100000; // [ 0.4453125]
storage[36] =  12'b010100100000; // [ 0.3203125]
storage[37] =  12'b010001110000; // [ 0.27734375]
storage[38] =  12'b010000110000; // [ 0.26171875]
storage[39] =  12'b010001110000; // [ 0.27734375]
storage[40] =  12'b010001110000; // [ 0.27734375]
storage[41] =  12'b010001110000; // [ 0.27734375]
storage[42] =  12'b010001110000; // [ 0.27734375]
storage[43] =  12'b010101000000; // [ 0.328125]
storage[44] =  12'b011101100000; // [ 0.4609375]
storage[45] =  12'b100101110000; // [ 0.58984375]
storage[46] =  12'b101000100000; // [ 0.6328125]
storage[47] =  12'b101001010000; // [ 0.64453125]
storage[48] =  12'b101001010000; // [ 0.64453125]
storage[49] =  12'b101001000000; // [ 0.640625]
storage[50] =  12'b101001010000; // [ 0.64453125]
storage[51] =  12'b101000110000; // [ 0.63671875]
storage[52] =  12'b101000110000; // [ 0.63671875]
storage[53] =  12'b101000010000; // [ 0.62890625]
storage[54] =  12'b101000000000; // [ 0.625]
storage[55] =  12'b100111100000; // [ 0.6171875]
storage[56] =  12'b100111000000; // [ 0.609375]
storage[57] =  12'b100111100000; // [ 0.6171875]
storage[58] =  12'b101000000000; // [ 0.625]
storage[59] =  12'b101000010000; // [ 0.62890625]
storage[60] =  12'b101000000000; // [ 0.625]
storage[61] =  12'b100110010000; // [ 0.59765625]
storage[62] =  12'b011101110000; // [ 0.46484375]
storage[63] =  12'b010010100000; // [ 0.2890625]
storage[64] =  12'b001111110000; // [ 0.24609375]
storage[65] =  12'b010100000000; // [ 0.3125]
storage[66] =  12'b011011010000; // [ 0.42578125]
storage[67] =  12'b011110110000; // [ 0.48046875]
storage[68] =  12'b011100010000; // [ 0.44140625]
storage[69] =  12'b010110010000; // [ 0.34765625]
storage[70] =  12'b010010000000; // [ 0.28125]
storage[71] =  12'b010000110000; // [ 0.26171875]
storage[72] =  12'b010101100000; // [ 0.3359375]
storage[73] =  12'b011111110000; // [ 0.49609375]
storage[74] =  12'b100111000000; // [ 0.609375]
storage[75] =  12'b101000110000; // [ 0.63671875]
storage[76] =  12'b101001000000; // [ 0.640625]
storage[77] =  12'b101001010000; // [ 0.64453125]
storage[78] =  12'b101001000000; // [ 0.640625]
storage[79] =  12'b101000110000; // [ 0.63671875]
storage[80] =  12'b101000100000; // [ 0.6328125]
storage[81] =  12'b101000010000; // [ 0.62890625]
storage[82] =  12'b101000000000; // [ 0.625]
storage[83] =  12'b100111110000; // [ 0.62109375]
storage[84] =  12'b100111010000; // [ 0.61328125]
storage[85] =  12'b100111100000; // [ 0.6171875]
storage[86] =  12'b100111110000; // [ 0.62109375]
storage[87] =  12'b100111110000; // [ 0.62109375]
storage[88] =  12'b100110110000; // [ 0.60546875]
storage[89] =  12'b100001000000; // [ 0.515625]
storage[90] =  12'b010011110000; // [ 0.30859375]
storage[91] =  12'b001111110000; // [ 0.24609375]
storage[92] =  12'b010101010000; // [ 0.33203125]
storage[93] =  12'b100000010000; // [ 0.50390625]
storage[94] =  12'b100111000000; // [ 0.609375]
storage[95] =  12'b101000010000; // [ 0.62890625]
storage[96] =  12'b100111000000; // [ 0.609375]
storage[97] =  12'b100001110000; // [ 0.52734375]
storage[98] =  12'b011001000000; // [ 0.390625]
storage[99] =  12'b010010100000; // [ 0.2890625]
storage[100] =  12'b010010010000; // [ 0.28515625]
storage[101] =  12'b011010010000; // [ 0.41015625]
storage[102] =  12'b100100000000; // [ 0.5625]
storage[103] =  12'b101000000000; // [ 0.625]
storage[104] =  12'b101000110000; // [ 0.63671875]
storage[105] =  12'b101001010000; // [ 0.64453125]
storage[106] =  12'b101001000000; // [ 0.640625]
storage[107] =  12'b101001000000; // [ 0.640625]
storage[108] =  12'b101000100000; // [ 0.6328125]
storage[109] =  12'b101000010000; // [ 0.62890625]
storage[110] =  12'b101000000000; // [ 0.625]
storage[111] =  12'b100111110000; // [ 0.62109375]
storage[112] =  12'b100111010000; // [ 0.61328125]
storage[113] =  12'b100111010000; // [ 0.61328125]
storage[114] =  12'b100111100000; // [ 0.6171875]
storage[115] =  12'b100111010000; // [ 0.61328125]
storage[116] =  12'b100100000000; // [ 0.5625]
storage[117] =  12'b010111000000; // [ 0.359375]
storage[118] =  12'b010000000000; // [ 0.25]
storage[119] =  12'b010010110000; // [ 0.29296875]
storage[120] =  12'b011110110000; // [ 0.48046875]
storage[121] =  12'b100111100000; // [ 0.6171875]
storage[122] =  12'b101001010000; // [ 0.64453125]
storage[123] =  12'b101001110000; // [ 0.65234375]
storage[124] =  12'b101010000000; // [ 0.65625]
storage[125] =  12'b100111010000; // [ 0.61328125]
storage[126] =  12'b100000010000; // [ 0.50390625]
storage[127] =  12'b010110110000; // [ 0.35546875]
storage[128] =  12'b010010100000; // [ 0.2890625]
storage[129] =  12'b010101110000; // [ 0.33984375]
storage[130] =  12'b100000100000; // [ 0.5078125]
storage[131] =  12'b100111000000; // [ 0.609375]
storage[132] =  12'b101000100000; // [ 0.6328125]
storage[133] =  12'b101001000000; // [ 0.640625]
storage[134] =  12'b101001010000; // [ 0.64453125]
storage[135] =  12'b101001000000; // [ 0.640625]
storage[136] =  12'b101000110000; // [ 0.63671875]
storage[137] =  12'b101000100000; // [ 0.6328125]
storage[138] =  12'b101000000000; // [ 0.625]
storage[139] =  12'b100111110000; // [ 0.62109375]
storage[140] =  12'b100111010000; // [ 0.61328125]
storage[141] =  12'b100111100000; // [ 0.6171875]
storage[142] =  12'b100111010000; // [ 0.61328125]
storage[143] =  12'b100110000000; // [ 0.59375]
storage[144] =  12'b011110010000; // [ 0.47265625]
storage[145] =  12'b010001110000; // [ 0.27734375]
storage[146] =  12'b010001100000; // [ 0.2734375]
storage[147] =  12'b011011000000; // [ 0.421875]
storage[148] =  12'b100101110000; // [ 0.58984375]
storage[149] =  12'b101000110000; // [ 0.63671875]
storage[150] =  12'b101010000000; // [ 0.65625]
storage[151] =  12'b101011000000; // [ 0.671875]
storage[152] =  12'b101010100000; // [ 0.6640625]
storage[153] =  12'b101010000000; // [ 0.65625]
storage[154] =  12'b100110010000; // [ 0.59765625]
storage[155] =  12'b011110110000; // [ 0.48046875]
storage[156] =  12'b010110010000; // [ 0.34765625]
storage[157] =  12'b010100110000; // [ 0.32421875]
storage[158] =  12'b011101010000; // [ 0.45703125]
storage[159] =  12'b100110000000; // [ 0.59375]
storage[160] =  12'b101000110000; // [ 0.63671875]
storage[161] =  12'b101001100000; // [ 0.6484375]
storage[162] =  12'b101001100000; // [ 0.6484375]
storage[163] =  12'b101001100000; // [ 0.6484375]
storage[164] =  12'b101001010000; // [ 0.64453125]
storage[165] =  12'b101000110000; // [ 0.63671875]
storage[166] =  12'b101000010000; // [ 0.62890625]
storage[167] =  12'b100111110000; // [ 0.62109375]
storage[168] =  12'b100111010000; // [ 0.61328125]
storage[169] =  12'b100111010000; // [ 0.61328125]
storage[170] =  12'b100111000000; // [ 0.609375]
storage[171] =  12'b100011110000; // [ 0.55859375]
storage[172] =  12'b010111100000; // [ 0.3671875]
storage[173] =  12'b010010000000; // [ 0.28125]
storage[174] =  12'b011000100000; // [ 0.3828125]
storage[175] =  12'b100100000000; // [ 0.5625]
storage[176] =  12'b101000100000; // [ 0.6328125]
storage[177] =  12'b101001110000; // [ 0.65234375]
storage[178] =  12'b101011000000; // [ 0.671875]
storage[179] =  12'b101011010000; // [ 0.67578125]
storage[180] =  12'b101011000000; // [ 0.671875]
storage[181] =  12'b101010110000; // [ 0.66796875]
storage[182] =  12'b101001110000; // [ 0.65234375]
storage[183] =  12'b100101000000; // [ 0.578125]
storage[184] =  12'b011100010000; // [ 0.44140625]
storage[185] =  12'b010101110000; // [ 0.33984375]
storage[186] =  12'b011011010000; // [ 0.42578125]
storage[187] =  12'b100100110000; // [ 0.57421875]
storage[188] =  12'b101000100000; // [ 0.6328125]
storage[189] =  12'b101010000000; // [ 0.65625]
storage[190] =  12'b101010000000; // [ 0.65625]
storage[191] =  12'b101010000000; // [ 0.65625]
storage[192] =  12'b101001100000; // [ 0.6484375]
storage[193] =  12'b101001000000; // [ 0.640625]
storage[194] =  12'b101000100000; // [ 0.6328125]
storage[195] =  12'b100111110000; // [ 0.62109375]
storage[196] =  12'b100111010000; // [ 0.61328125]
storage[197] =  12'b100111100000; // [ 0.6171875]
storage[198] =  12'b100110010000; // [ 0.59765625]
storage[199] =  12'b011111110000; // [ 0.49609375]
storage[200] =  12'b010011100000; // [ 0.3046875]
storage[201] =  12'b010100000000; // [ 0.3125]
storage[202] =  12'b011110110000; // [ 0.48046875]
storage[203] =  12'b100111110000; // [ 0.62109375]
storage[204] =  12'b101001100000; // [ 0.6484375]
storage[205] =  12'b101010110000; // [ 0.66796875]
storage[206] =  12'b101011110000; // [ 0.68359375]
storage[207] =  12'b101011110000; // [ 0.68359375]
storage[208] =  12'b101011100000; // [ 0.6796875]
storage[209] =  12'b101011010000; // [ 0.67578125]
storage[210] =  12'b101010110000; // [ 0.66796875]
storage[211] =  12'b101000000000; // [ 0.625]
storage[212] =  12'b100000000000; // [ 0.5]
storage[213] =  12'b010111010000; // [ 0.36328125]
storage[214] =  12'b011010100000; // [ 0.4140625]
storage[215] =  12'b100100000000; // [ 0.5625]
storage[216] =  12'b101000100000; // [ 0.6328125]
storage[217] =  12'b101010000000; // [ 0.65625]
storage[218] =  12'b101010100000; // [ 0.6640625]
storage[219] =  12'b101010000000; // [ 0.65625]
storage[220] =  12'b101010000000; // [ 0.65625]
storage[221] =  12'b101001000000; // [ 0.640625]
storage[222] =  12'b101000110000; // [ 0.63671875]
storage[223] =  12'b101000000000; // [ 0.625]
storage[224] =  12'b100111100000; // [ 0.6171875]
storage[225] =  12'b100111010000; // [ 0.61328125]
storage[226] =  12'b100101010000; // [ 0.58203125]
storage[227] =  12'b011011010000; // [ 0.42578125]
storage[228] =  12'b010010000000; // [ 0.28125]
storage[229] =  12'b010111010000; // [ 0.36328125]
storage[230] =  12'b100011010000; // [ 0.55078125]
storage[231] =  12'b101000110000; // [ 0.63671875]
storage[232] =  12'b101010110000; // [ 0.66796875]
storage[233] =  12'b101011100000; // [ 0.6796875]
storage[234] =  12'b101100000000; // [ 0.6875]
storage[235] =  12'b101100000000; // [ 0.6875]
storage[236] =  12'b101100000000; // [ 0.6875]
storage[237] =  12'b101011110000; // [ 0.68359375]
storage[238] =  12'b101011000000; // [ 0.671875]
storage[239] =  12'b101001010000; // [ 0.64453125]
storage[240] =  12'b100010000000; // [ 0.53125]
storage[241] =  12'b011000100000; // [ 0.3828125]
storage[242] =  12'b011001010000; // [ 0.39453125]
storage[243] =  12'b100011000000; // [ 0.546875]
storage[244] =  12'b101000010000; // [ 0.62890625]
storage[245] =  12'b101010010000; // [ 0.66015625]
storage[246] =  12'b101010100000; // [ 0.6640625]
storage[247] =  12'b101010110000; // [ 0.66796875]
storage[248] =  12'b101001110000; // [ 0.65234375]
storage[249] =  12'b101001100000; // [ 0.6484375]
storage[250] =  12'b101000110000; // [ 0.63671875]
storage[251] =  12'b101000000000; // [ 0.625]
storage[252] =  12'b100111000000; // [ 0.609375]
storage[253] =  12'b100111000000; // [ 0.609375]
storage[254] =  12'b100011110000; // [ 0.55859375]
storage[255] =  12'b010111110000; // [ 0.37109375]
storage[256] =  12'b010010000000; // [ 0.28125]
storage[257] =  12'b011011010000; // [ 0.42578125]
storage[258] =  12'b100110110000; // [ 0.60546875]
storage[259] =  12'b101001110000; // [ 0.65234375]
storage[260] =  12'b101011010000; // [ 0.67578125]
storage[261] =  12'b101100000000; // [ 0.6875]
storage[262] =  12'b101100000000; // [ 0.6875]
storage[263] =  12'b101100000000; // [ 0.6875]
storage[264] =  12'b101100000000; // [ 0.6875]
storage[265] =  12'b101100000000; // [ 0.6875]
storage[266] =  12'b101011100000; // [ 0.6796875]
storage[267] =  12'b101010000000; // [ 0.65625]
storage[268] =  12'b100011000000; // [ 0.546875]
storage[269] =  12'b011001100000; // [ 0.3984375]
storage[270] =  12'b010111000000; // [ 0.359375]
storage[271] =  12'b100001100000; // [ 0.5234375]
storage[272] =  12'b100111110000; // [ 0.62109375]
storage[273] =  12'b101010000000; // [ 0.65625]
storage[274] =  12'b101010100000; // [ 0.6640625]
storage[275] =  12'b101010010000; // [ 0.66015625]
storage[276] =  12'b101010000000; // [ 0.65625]
storage[277] =  12'b101001100000; // [ 0.6484375]
storage[278] =  12'b101000100000; // [ 0.6328125]
storage[279] =  12'b101000010000; // [ 0.62890625]
storage[280] =  12'b100111000000; // [ 0.609375]
storage[281] =  12'b100110100000; // [ 0.6015625]
storage[282] =  12'b100001100000; // [ 0.5234375]
storage[283] =  12'b010100110000; // [ 0.32421875]
storage[284] =  12'b010011010000; // [ 0.30078125]
storage[285] =  12'b011110100000; // [ 0.4765625]
storage[286] =  12'b101000000000; // [ 0.625]
storage[287] =  12'b101010000000; // [ 0.65625]
storage[288] =  12'b101011100000; // [ 0.6796875]
storage[289] =  12'b101011110000; // [ 0.68359375]
storage[290] =  12'b101100000000; // [ 0.6875]
storage[291] =  12'b101100000000; // [ 0.6875]
storage[292] =  12'b101100010000; // [ 0.69140625]
storage[293] =  12'b101100000000; // [ 0.6875]
storage[294] =  12'b101011100000; // [ 0.6796875]
storage[295] =  12'b101010010000; // [ 0.66015625]
storage[296] =  12'b100011110000; // [ 0.55859375]
storage[297] =  12'b011010000000; // [ 0.40625]
storage[298] =  12'b010101110000; // [ 0.33984375]
storage[299] =  12'b100000100000; // [ 0.5078125]
storage[300] =  12'b100111100000; // [ 0.6171875]
storage[301] =  12'b101001110000; // [ 0.65234375]
storage[302] =  12'b101010100000; // [ 0.6640625]
storage[303] =  12'b101010010000; // [ 0.66015625]
storage[304] =  12'b101001110000; // [ 0.65234375]
storage[305] =  12'b101001100000; // [ 0.6484375]
storage[306] =  12'b101000100000; // [ 0.6328125]
storage[307] =  12'b101000000000; // [ 0.625]
storage[308] =  12'b100111010000; // [ 0.61328125]
storage[309] =  12'b100110000000; // [ 0.59375]
storage[310] =  12'b011111000000; // [ 0.484375]
storage[311] =  12'b010011000000; // [ 0.296875]
storage[312] =  12'b010100110000; // [ 0.32421875]
storage[313] =  12'b100010010000; // [ 0.53515625]
storage[314] =  12'b101000100000; // [ 0.6328125]
storage[315] =  12'b101010100000; // [ 0.6640625]
storage[316] =  12'b101011010000; // [ 0.67578125]
storage[317] =  12'b101011100000; // [ 0.6796875]
storage[318] =  12'b101011100000; // [ 0.6796875]
storage[319] =  12'b101100000000; // [ 0.6875]
storage[320] =  12'b101100000000; // [ 0.6875]
storage[321] =  12'b101100000000; // [ 0.6875]
storage[322] =  12'b101011100000; // [ 0.6796875]
storage[323] =  12'b101010010000; // [ 0.66015625]
storage[324] =  12'b100011100000; // [ 0.5546875]
storage[325] =  12'b011010000000; // [ 0.40625]
storage[326] =  12'b010101100000; // [ 0.3359375]
storage[327] =  12'b100000000000; // [ 0.5]
storage[328] =  12'b100111010000; // [ 0.61328125]
storage[329] =  12'b101001100000; // [ 0.6484375]
storage[330] =  12'b101010000000; // [ 0.65625]
storage[331] =  12'b101010000000; // [ 0.65625]
storage[332] =  12'b101001110000; // [ 0.65234375]
storage[333] =  12'b101001000000; // [ 0.640625]
storage[334] =  12'b101000010000; // [ 0.62890625]
storage[335] =  12'b100111110000; // [ 0.62109375]
storage[336] =  12'b100111000000; // [ 0.609375]
storage[337] =  12'b100101000000; // [ 0.578125]
storage[338] =  12'b011011110000; // [ 0.43359375]
storage[339] =  12'b010001110000; // [ 0.27734375]
storage[340] =  12'b010111000000; // [ 0.359375]
storage[341] =  12'b100011110000; // [ 0.55859375]
storage[342] =  12'b101001000000; // [ 0.640625]
storage[343] =  12'b101010010000; // [ 0.66015625]
storage[344] =  12'b101011000000; // [ 0.671875]
storage[345] =  12'b101011000000; // [ 0.671875]
storage[346] =  12'b101011010000; // [ 0.67578125]
storage[347] =  12'b101011100000; // [ 0.6796875]
storage[348] =  12'b101011100000; // [ 0.6796875]
storage[349] =  12'b101011100000; // [ 0.6796875]
storage[350] =  12'b101010110000; // [ 0.66796875]
storage[351] =  12'b101001100000; // [ 0.6484375]
storage[352] =  12'b100011010000; // [ 0.55078125]
storage[353] =  12'b011001100000; // [ 0.3984375]
storage[354] =  12'b010101010000; // [ 0.33203125]
storage[355] =  12'b100000100000; // [ 0.5078125]
storage[356] =  12'b100111010000; // [ 0.61328125]
storage[357] =  12'b101001000000; // [ 0.640625]
storage[358] =  12'b101010000000; // [ 0.65625]
storage[359] =  12'b101001110000; // [ 0.65234375]
storage[360] =  12'b101001010000; // [ 0.64453125]
storage[361] =  12'b101000110000; // [ 0.63671875]
storage[362] =  12'b101000010000; // [ 0.62890625]
storage[363] =  12'b100111100000; // [ 0.6171875]
storage[364] =  12'b100110100000; // [ 0.6015625]
storage[365] =  12'b100100000000; // [ 0.5625]
storage[366] =  12'b011001000000; // [ 0.390625]
storage[367] =  12'b010001110000; // [ 0.27734375]
storage[368] =  12'b011001100000; // [ 0.3984375]
storage[369] =  12'b100101010000; // [ 0.58203125]
storage[370] =  12'b101000110000; // [ 0.63671875]
storage[371] =  12'b101010000000; // [ 0.65625]
storage[372] =  12'b101010110000; // [ 0.66796875]
storage[373] =  12'b101010110000; // [ 0.66796875]
storage[374] =  12'b101010110000; // [ 0.66796875]
storage[375] =  12'b101011000000; // [ 0.671875]
storage[376] =  12'b101011010000; // [ 0.67578125]
storage[377] =  12'b101010110000; // [ 0.66796875]
storage[378] =  12'b101010010000; // [ 0.66015625]
storage[379] =  12'b101000110000; // [ 0.63671875]
storage[380] =  12'b100010100000; // [ 0.5390625]
storage[381] =  12'b011000100000; // [ 0.3828125]
storage[382] =  12'b010101110000; // [ 0.33984375]
storage[383] =  12'b100001100000; // [ 0.5234375]
storage[384] =  12'b100111100000; // [ 0.6171875]
storage[385] =  12'b101001010000; // [ 0.64453125]
storage[386] =  12'b101001010000; // [ 0.64453125]
storage[387] =  12'b101001010000; // [ 0.64453125]
storage[388] =  12'b101001000000; // [ 0.640625]
storage[389] =  12'b101000100000; // [ 0.6328125]
storage[390] =  12'b101000000000; // [ 0.625]
storage[391] =  12'b100111100000; // [ 0.6171875]
storage[392] =  12'b100110010000; // [ 0.59765625]
storage[393] =  12'b100011000000; // [ 0.546875]
storage[394] =  12'b010111110000; // [ 0.37109375]
storage[395] =  12'b010001110000; // [ 0.27734375]
storage[396] =  12'b011011000000; // [ 0.421875]
storage[397] =  12'b100110000000; // [ 0.59375]
storage[398] =  12'b101001000000; // [ 0.640625]
storage[399] =  12'b101001110000; // [ 0.65234375]
storage[400] =  12'b101010010000; // [ 0.66015625]
storage[401] =  12'b101010100000; // [ 0.6640625]
storage[402] =  12'b101011000000; // [ 0.671875]
storage[403] =  12'b101011000000; // [ 0.671875]
storage[404] =  12'b101011000000; // [ 0.671875]
storage[405] =  12'b101010110000; // [ 0.66796875]
storage[406] =  12'b101010010000; // [ 0.66015625]
storage[407] =  12'b100111110000; // [ 0.62109375]
storage[408] =  12'b100000000000; // [ 0.5]
storage[409] =  12'b010101110000; // [ 0.33984375]
storage[410] =  12'b010110100000; // [ 0.3515625]
storage[411] =  12'b100010100000; // [ 0.5390625]
storage[412] =  12'b100111110000; // [ 0.62109375]
storage[413] =  12'b101001010000; // [ 0.64453125]
storage[414] =  12'b101001010000; // [ 0.64453125]
storage[415] =  12'b101001010000; // [ 0.64453125]
storage[416] =  12'b101000110000; // [ 0.63671875]
storage[417] =  12'b101000010000; // [ 0.62890625]
storage[418] =  12'b100111110000; // [ 0.62109375]
storage[419] =  12'b100111010000; // [ 0.61328125]
storage[420] =  12'b100110010000; // [ 0.59765625]
storage[421] =  12'b100010100000; // [ 0.5390625]
storage[422] =  12'b010111110000; // [ 0.37109375]
storage[423] =  12'b010010100000; // [ 0.2890625]
storage[424] =  12'b011011010000; // [ 0.42578125]
storage[425] =  12'b100110010000; // [ 0.59765625]
storage[426] =  12'b101000110000; // [ 0.63671875]
storage[427] =  12'b101001110000; // [ 0.65234375]
storage[428] =  12'b101010000000; // [ 0.65625]
storage[429] =  12'b101010010000; // [ 0.66015625]
storage[430] =  12'b101010100000; // [ 0.6640625]
storage[431] =  12'b101010100000; // [ 0.6640625]
storage[432] =  12'b101010110000; // [ 0.66796875]
storage[433] =  12'b101010110000; // [ 0.66796875]
storage[434] =  12'b101010010000; // [ 0.66015625]
storage[435] =  12'b100110100000; // [ 0.6015625]
storage[436] =  12'b011101000000; // [ 0.453125]
storage[437] =  12'b010011000000; // [ 0.296875]
storage[438] =  12'b010111000000; // [ 0.359375]
storage[439] =  12'b100011010000; // [ 0.55078125]
storage[440] =  12'b101000000000; // [ 0.625]
storage[441] =  12'b101001000000; // [ 0.640625]
storage[442] =  12'b101001000000; // [ 0.640625]
storage[443] =  12'b101001000000; // [ 0.640625]
storage[444] =  12'b101000100000; // [ 0.6328125]
storage[445] =  12'b101000000000; // [ 0.625]
storage[446] =  12'b100111100000; // [ 0.6171875]
storage[447] =  12'b100111010000; // [ 0.61328125]
storage[448] =  12'b100110000000; // [ 0.59375]
storage[449] =  12'b100011000000; // [ 0.546875]
storage[450] =  12'b011001000000; // [ 0.390625]
storage[451] =  12'b010010100000; // [ 0.2890625]
storage[452] =  12'b011010010000; // [ 0.41015625]
storage[453] =  12'b100101000000; // [ 0.578125]
storage[454] =  12'b101000100000; // [ 0.6328125]
storage[455] =  12'b101001000000; // [ 0.640625]
storage[456] =  12'b101001110000; // [ 0.65234375]
storage[457] =  12'b101001100000; // [ 0.6484375]
storage[458] =  12'b101001110000; // [ 0.65234375]
storage[459] =  12'b101010100000; // [ 0.6640625]
storage[460] =  12'b101010100000; // [ 0.6640625]
storage[461] =  12'b101010100000; // [ 0.6640625]
storage[462] =  12'b101001110000; // [ 0.65234375]
storage[463] =  12'b100011110000; // [ 0.55859375]
storage[464] =  12'b011000100000; // [ 0.3828125]
storage[465] =  12'b010001100000; // [ 0.2734375]
storage[466] =  12'b011000100000; // [ 0.3828125]
storage[467] =  12'b100100000000; // [ 0.5625]
storage[468] =  12'b101000000000; // [ 0.625]
storage[469] =  12'b101000110000; // [ 0.63671875]
storage[470] =  12'b101000110000; // [ 0.63671875]
storage[471] =  12'b101000100000; // [ 0.6328125]
storage[472] =  12'b101000000000; // [ 0.625]
storage[473] =  12'b100111110000; // [ 0.62109375]
storage[474] =  12'b100111100000; // [ 0.6171875]
storage[475] =  12'b100111000000; // [ 0.609375]
storage[476] =  12'b100110100000; // [ 0.6015625]
storage[477] =  12'b100100010000; // [ 0.56640625]
storage[478] =  12'b011100010000; // [ 0.44140625]
storage[479] =  12'b010011000000; // [ 0.296875]
storage[480] =  12'b011001100000; // [ 0.3984375]
storage[481] =  12'b100100100000; // [ 0.5703125]
storage[482] =  12'b101000000000; // [ 0.625]
storage[483] =  12'b101001010000; // [ 0.64453125]
storage[484] =  12'b101001010000; // [ 0.64453125]
storage[485] =  12'b101001110000; // [ 0.65234375]
storage[486] =  12'b101010000000; // [ 0.65625]
storage[487] =  12'b101010100000; // [ 0.6640625]
storage[488] =  12'b101010110000; // [ 0.66796875]
storage[489] =  12'b101010010000; // [ 0.66015625]
storage[490] =  12'b100111100000; // [ 0.6171875]
storage[491] =  12'b011110010000; // [ 0.47265625]
storage[492] =  12'b010011010000; // [ 0.30078125]
storage[493] =  12'b010001000000; // [ 0.265625]
storage[494] =  12'b011100100000; // [ 0.4453125]
storage[495] =  12'b100110000000; // [ 0.59375]
storage[496] =  12'b101000110000; // [ 0.63671875]
storage[497] =  12'b101001000000; // [ 0.640625]
storage[498] =  12'b101001010000; // [ 0.64453125]
storage[499] =  12'b101000110000; // [ 0.63671875]
storage[500] =  12'b101000010000; // [ 0.62890625]
storage[501] =  12'b100111110000; // [ 0.62109375]
storage[502] =  12'b100111100000; // [ 0.6171875]
storage[503] =  12'b100111010000; // [ 0.61328125]
storage[504] =  12'b100110110000; // [ 0.60546875]
storage[505] =  12'b100101000000; // [ 0.578125]
storage[506] =  12'b011111010000; // [ 0.48828125]
storage[507] =  12'b010100100000; // [ 0.3203125]
storage[508] =  12'b011000100000; // [ 0.3828125]
storage[509] =  12'b100011100000; // [ 0.5546875]
storage[510] =  12'b100111110000; // [ 0.62109375]
storage[511] =  12'b101000110000; // [ 0.63671875]
storage[512] =  12'b101001010000; // [ 0.64453125]
storage[513] =  12'b101001100000; // [ 0.6484375]
storage[514] =  12'b101010000000; // [ 0.65625]
storage[515] =  12'b101010100000; // [ 0.6640625]
storage[516] =  12'b101010100000; // [ 0.6640625]
storage[517] =  12'b101010000000; // [ 0.65625]
storage[518] =  12'b100011010000; // [ 0.55078125]
storage[519] =  12'b010111110000; // [ 0.37109375]
storage[520] =  12'b010000000000; // [ 0.25]
storage[521] =  12'b010010000000; // [ 0.28125]
storage[522] =  12'b100000110000; // [ 0.51171875]
storage[523] =  12'b100111010000; // [ 0.61328125]
storage[524] =  12'b101001000000; // [ 0.640625]
storage[525] =  12'b101001100000; // [ 0.6484375]
storage[526] =  12'b101000110000; // [ 0.63671875]
storage[527] =  12'b101000110000; // [ 0.63671875]
storage[528] =  12'b101000010000; // [ 0.62890625]
storage[529] =  12'b100111110000; // [ 0.62109375]
storage[530] =  12'b100111100000; // [ 0.6171875]
storage[531] =  12'b100111000000; // [ 0.609375]
storage[532] =  12'b100110010000; // [ 0.59765625]
storage[533] =  12'b100101010000; // [ 0.58203125]
storage[534] =  12'b100001100000; // [ 0.5234375]
storage[535] =  12'b010111100000; // [ 0.3671875]
storage[536] =  12'b010101110000; // [ 0.33984375]
storage[537] =  12'b100000100000; // [ 0.5078125]
storage[538] =  12'b100111000000; // [ 0.609375]
storage[539] =  12'b101000010000; // [ 0.62890625]
storage[540] =  12'b101000110000; // [ 0.63671875]
storage[541] =  12'b101001010000; // [ 0.64453125]
storage[542] =  12'b101001100000; // [ 0.6484375]
storage[543] =  12'b101010010000; // [ 0.66015625]
storage[544] =  12'b101010010000; // [ 0.66015625]
storage[545] =  12'b100111110000; // [ 0.62109375]
storage[546] =  12'b011111000000; // [ 0.484375]
storage[547] =  12'b010010110000; // [ 0.29296875]
storage[548] =  12'b001110100000; // [ 0.2265625]
storage[549] =  12'b010100100000; // [ 0.3203125]
storage[550] =  12'b100010110000; // [ 0.54296875]
storage[551] =  12'b100111110000; // [ 0.62109375]
storage[552] =  12'b101001010000; // [ 0.64453125]
storage[553] =  12'b101000110000; // [ 0.63671875]
storage[554] =  12'b101000100000; // [ 0.6328125]
storage[555] =  12'b101000000000; // [ 0.625]
storage[556] =  12'b100111100000; // [ 0.6171875]
storage[557] =  12'b100111010000; // [ 0.61328125]
storage[558] =  12'b100111000000; // [ 0.609375]
storage[559] =  12'b100110110000; // [ 0.60546875]
storage[560] =  12'b100101110000; // [ 0.58984375]
storage[561] =  12'b100101100000; // [ 0.5859375]
storage[562] =  12'b100011010000; // [ 0.55078125]
storage[563] =  12'b011011110000; // [ 0.43359375]
storage[564] =  12'b010101000000; // [ 0.328125]
storage[565] =  12'b011100100000; // [ 0.4453125]
storage[566] =  12'b100101110000; // [ 0.58984375]
storage[567] =  12'b100111110000; // [ 0.62109375]
storage[568] =  12'b101000100000; // [ 0.6328125]
storage[569] =  12'b101000110000; // [ 0.63671875]
storage[570] =  12'b101001110000; // [ 0.65234375]
storage[571] =  12'b101001110000; // [ 0.65234375]
storage[572] =  12'b101010000000; // [ 0.65625]
storage[573] =  12'b100101110000; // [ 0.58984375]
storage[574] =  12'b011011010000; // [ 0.42578125]
storage[575] =  12'b010000100000; // [ 0.2578125]
storage[576] =  12'b001110100000; // [ 0.2265625]
storage[577] =  12'b011000010000; // [ 0.37890625]
storage[578] =  12'b100100110000; // [ 0.57421875]
storage[579] =  12'b101000010000; // [ 0.62890625]
storage[580] =  12'b101001010000; // [ 0.64453125]
storage[581] =  12'b101000100000; // [ 0.6328125]
storage[582] =  12'b101000000000; // [ 0.625]
storage[583] =  12'b100111110000; // [ 0.62109375]
storage[584] =  12'b100111100000; // [ 0.6171875]
storage[585] =  12'b100111000000; // [ 0.609375]
storage[586] =  12'b100110100000; // [ 0.6015625]
storage[587] =  12'b100110010000; // [ 0.59765625]
storage[588] =  12'b100101110000; // [ 0.58984375]
storage[589] =  12'b100101110000; // [ 0.58984375]
storage[590] =  12'b100100110000; // [ 0.57421875]
storage[591] =  12'b100000100000; // [ 0.5078125]
storage[592] =  12'b010111000000; // [ 0.359375]
storage[593] =  12'b011000110000; // [ 0.38671875]
storage[594] =  12'b100010100000; // [ 0.5390625]
storage[595] =  12'b100111010000; // [ 0.61328125]
storage[596] =  12'b101000010000; // [ 0.62890625]
storage[597] =  12'b101000110000; // [ 0.63671875]
storage[598] =  12'b101001000000; // [ 0.640625]
storage[599] =  12'b101001010000; // [ 0.64453125]
storage[600] =  12'b100111110000; // [ 0.62109375]
storage[601] =  12'b100000000000; // [ 0.5]
storage[602] =  12'b010100100000; // [ 0.3203125]
storage[603] =  12'b001110010000; // [ 0.22265625]
storage[604] =  12'b010000000000; // [ 0.25]
storage[605] =  12'b011101100000; // [ 0.4609375]
storage[606] =  12'b100110100000; // [ 0.6015625]
storage[607] =  12'b101000100000; // [ 0.6328125]
storage[608] =  12'b101000110000; // [ 0.63671875]
storage[609] =  12'b101000010000; // [ 0.62890625]
storage[610] =  12'b101000000000; // [ 0.625]
storage[611] =  12'b100111110000; // [ 0.62109375]
storage[612] =  12'b100111010000; // [ 0.61328125]
storage[613] =  12'b100110110000; // [ 0.60546875]
storage[614] =  12'b100110010000; // [ 0.59765625]
storage[615] =  12'b100101110000; // [ 0.58984375]
storage[616] =  12'b100101100000; // [ 0.5859375]
storage[617] =  12'b100101100000; // [ 0.5859375]
storage[618] =  12'b100101100000; // [ 0.5859375]
storage[619] =  12'b100011010000; // [ 0.55078125]
storage[620] =  12'b011100110000; // [ 0.44921875]
storage[621] =  12'b010101010000; // [ 0.33203125]
storage[622] =  12'b011011100000; // [ 0.4296875]
storage[623] =  12'b100100000000; // [ 0.5625]
storage[624] =  12'b100111000000; // [ 0.609375]
storage[625] =  12'b101000000000; // [ 0.625]
storage[626] =  12'b101000000000; // [ 0.625]
storage[627] =  12'b100111100000; // [ 0.6171875]
storage[628] =  12'b100010000000; // [ 0.53125]
storage[629] =  12'b010110010000; // [ 0.34765625]
storage[630] =  12'b001110100000; // [ 0.2265625]
storage[631] =  12'b001110100000; // [ 0.2265625]
storage[632] =  12'b010101010000; // [ 0.33203125]
storage[633] =  12'b100010000000; // [ 0.53125]
storage[634] =  12'b100111000000; // [ 0.609375]
storage[635] =  12'b101000000000; // [ 0.625]
storage[636] =  12'b101000000000; // [ 0.625]
storage[637] =  12'b100111110000; // [ 0.62109375]
storage[638] =  12'b100111010000; // [ 0.61328125]
storage[639] =  12'b100111000000; // [ 0.609375]
storage[640] =  12'b100110100000; // [ 0.6015625]
storage[641] =  12'b100101110000; // [ 0.58984375]
storage[642] =  12'b100101100000; // [ 0.5859375]
storage[643] =  12'b100101010000; // [ 0.58203125]
storage[644] =  12'b100101000000; // [ 0.578125]
storage[645] =  12'b100101000000; // [ 0.578125]
storage[646] =  12'b100101100000; // [ 0.5859375]
storage[647] =  12'b100100110000; // [ 0.57421875]
storage[648] =  12'b100001000000; // [ 0.515625]
storage[649] =  12'b010111000000; // [ 0.359375]
storage[650] =  12'b010011000000; // [ 0.296875]
storage[651] =  12'b011000000000; // [ 0.375]
storage[652] =  12'b011111100000; // [ 0.4921875]
storage[653] =  12'b100100010000; // [ 0.56640625]
storage[654] =  12'b100100110000; // [ 0.57421875]
storage[655] =  12'b100001000000; // [ 0.515625]
storage[656] =  12'b010111110000; // [ 0.37109375]
storage[657] =  12'b001111100000; // [ 0.2421875]
storage[658] =  12'b001110010000; // [ 0.22265625]
storage[659] =  12'b010011010000; // [ 0.30078125]
storage[660] =  12'b011110100000; // [ 0.4765625]
storage[661] =  12'b100110000000; // [ 0.59375]
storage[662] =  12'b100111100000; // [ 0.6171875]
storage[663] =  12'b100111100000; // [ 0.6171875]
storage[664] =  12'b100111100000; // [ 0.6171875]
storage[665] =  12'b100111010000; // [ 0.61328125]
storage[666] =  12'b100111000000; // [ 0.609375]
storage[667] =  12'b100110100000; // [ 0.6015625]
storage[668] =  12'b100110000000; // [ 0.59375]
storage[669] =  12'b100101110000; // [ 0.58984375]
storage[670] =  12'b100101100000; // [ 0.5859375]
storage[671] =  12'b100100110000; // [ 0.57421875]
storage[672] =  12'b100100110000; // [ 0.57421875]
storage[673] =  12'b100101010000; // [ 0.58203125]
storage[674] =  12'b100101100000; // [ 0.5859375]
storage[675] =  12'b100101100000; // [ 0.5859375]
storage[676] =  12'b100011110000; // [ 0.55859375]
storage[677] =  12'b011101110000; // [ 0.46484375]
storage[678] =  12'b010010110000; // [ 0.29296875]
storage[679] =  12'b001111010000; // [ 0.23828125]
storage[680] =  12'b010010000000; // [ 0.28125]
storage[681] =  12'b010101000000; // [ 0.328125]
storage[682] =  12'b010101010000; // [ 0.33203125]
storage[683] =  12'b010010000000; // [ 0.28125]
storage[684] =  12'b001111000000; // [ 0.234375]
storage[685] =  12'b001111010000; // [ 0.23828125]
storage[686] =  12'b010100100000; // [ 0.3203125]
storage[687] =  12'b011110100000; // [ 0.4765625]
storage[688] =  12'b100101110000; // [ 0.58984375]
storage[689] =  12'b100111010000; // [ 0.61328125]
storage[690] =  12'b100111100000; // [ 0.6171875]
storage[691] =  12'b100111000000; // [ 0.609375]
storage[692] =  12'b100111010000; // [ 0.61328125]
storage[693] =  12'b100111000000; // [ 0.609375]
storage[694] =  12'b100110100000; // [ 0.6015625]
storage[695] =  12'b100110010000; // [ 0.59765625]
storage[696] =  12'b100101110000; // [ 0.58984375]
storage[697] =  12'b100101100000; // [ 0.5859375]
storage[698] =  12'b100101010000; // [ 0.58203125]
storage[699] =  12'b100100100000; // [ 0.5703125]
storage[700] =  12'b100100010000; // [ 0.56640625]
storage[701] =  12'b100100110000; // [ 0.57421875]
storage[702] =  12'b100101010000; // [ 0.58203125]
storage[703] =  12'b100101100000; // [ 0.5859375]
storage[704] =  12'b100101000000; // [ 0.578125]
storage[705] =  12'b100011000000; // [ 0.546875]
storage[706] =  12'b011100000000; // [ 0.4375]
storage[707] =  12'b010010000000; // [ 0.28125]
storage[708] =  12'b001101110000; // [ 0.21484375]
storage[709] =  12'b001101010000; // [ 0.20703125]
storage[710] =  12'b001101100000; // [ 0.2109375]
storage[711] =  12'b001111000000; // [ 0.234375]
storage[712] =  12'b010010000000; // [ 0.28125]
storage[713] =  12'b011001000000; // [ 0.390625]
storage[714] =  12'b100001000000; // [ 0.515625]
storage[715] =  12'b100110000000; // [ 0.59375]
storage[716] =  12'b100111000000; // [ 0.609375]
storage[717] =  12'b100111000000; // [ 0.609375]
storage[718] =  12'b100111000000; // [ 0.609375]
storage[719] =  12'b100110110000; // [ 0.60546875]
storage[720] =  12'b100110110000; // [ 0.60546875]
storage[721] =  12'b100110100000; // [ 0.6015625]
storage[722] =  12'b100110010000; // [ 0.59765625]
storage[723] =  12'b100101110000; // [ 0.58984375]
storage[724] =  12'b100101010000; // [ 0.58203125]
storage[725] =  12'b100101000000; // [ 0.578125]
storage[726] =  12'b100100110000; // [ 0.57421875]
storage[727] =  12'b100100000000; // [ 0.5625]
storage[728] =  12'b100011110000; // [ 0.55859375]
storage[729] =  12'b100100100000; // [ 0.5703125]
storage[730] =  12'b100100110000; // [ 0.57421875]
storage[731] =  12'b100101000000; // [ 0.578125]
storage[732] =  12'b100101010000; // [ 0.58203125]
storage[733] =  12'b100101000000; // [ 0.578125]
storage[734] =  12'b100011000000; // [ 0.546875]
storage[735] =  12'b011101110000; // [ 0.46484375]
storage[736] =  12'b010110100000; // [ 0.3515625]
storage[737] =  12'b010010100000; // [ 0.2890625]
storage[738] =  12'b010011110000; // [ 0.30859375]
storage[739] =  12'b011001010000; // [ 0.39453125]
storage[740] =  12'b100000010000; // [ 0.50390625]
storage[741] =  12'b100100110000; // [ 0.57421875]
storage[742] =  12'b100110110000; // [ 0.60546875]
storage[743] =  12'b100111000000; // [ 0.609375]
storage[744] =  12'b100110110000; // [ 0.60546875]
storage[745] =  12'b100110110000; // [ 0.60546875]
storage[746] =  12'b100110100000; // [ 0.6015625]
storage[747] =  12'b100110100000; // [ 0.6015625]
storage[748] =  12'b100110100000; // [ 0.6015625]
storage[749] =  12'b100110010000; // [ 0.59765625]
storage[750] =  12'b100101110000; // [ 0.58984375]
storage[751] =  12'b100101010000; // [ 0.58203125]
storage[752] =  12'b100101000000; // [ 0.578125]
storage[753] =  12'b100100110000; // [ 0.57421875]
storage[754] =  12'b100100010000; // [ 0.56640625]
storage[755] =  12'b100011100000; // [ 0.5546875]
storage[756] =  12'b100011010000; // [ 0.55078125]
storage[757] =  12'b100011110000; // [ 0.55859375]
storage[758] =  12'b100100100000; // [ 0.5703125]
storage[759] =  12'b100101000000; // [ 0.578125]
storage[760] =  12'b100101100000; // [ 0.5859375]
storage[761] =  12'b100101110000; // [ 0.58984375]
storage[762] =  12'b100110000000; // [ 0.59375]
storage[763] =  12'b100101000000; // [ 0.578125]
storage[764] =  12'b100011000000; // [ 0.546875]
storage[765] =  12'b100001100000; // [ 0.5234375]
storage[766] =  12'b100010100000; // [ 0.5390625]
storage[767] =  12'b100101000000; // [ 0.578125]
storage[768] =  12'b100110100000; // [ 0.6015625]
storage[769] =  12'b100111000000; // [ 0.609375]
storage[770] =  12'b100111000000; // [ 0.609375]
storage[771] =  12'b100110110000; // [ 0.60546875]
storage[772] =  12'b100110100000; // [ 0.6015625]
storage[773] =  12'b100110010000; // [ 0.59765625]
storage[774] =  12'b100110010000; // [ 0.59765625]
storage[775] =  12'b100110010000; // [ 0.59765625]
storage[776] =  12'b100110000000; // [ 0.59375]
storage[777] =  12'b100101110000; // [ 0.58984375]
storage[778] =  12'b100101010000; // [ 0.58203125]
storage[779] =  12'b100101000000; // [ 0.578125]
storage[780] =  12'b100100110000; // [ 0.57421875]
storage[781] =  12'b100100100000; // [ 0.5703125]
storage[782] =  12'b100100000000; // [ 0.5625]
storage[783] =  12'b100011010000; // [ 0.55078125]
storage[784] =  13'b0001100111011; // 827 0.20187625288963318
storage[785] =  13'b0100000010001; // 2065 0.504081130027771
storage[786] =  13'b0000010011001; // 153 0.037423789501190186
storage[787] =  13'b0000110111010; // 442 0.10783947259187698
storage[788] = -13'b0000100100011; // -291 -0.07114624232053757
storage[789] = -13'b0001111011000; // -984 -0.24016837775707245
storage[790] = -13'b0000011011100; // -220 -0.05364435166120529
storage[791] = -13'b0011001000101; // -1605 -0.391905277967453
storage[792] = -13'b0001001111110; // -638 -0.15579168498516083
storage[793] =  13'b0010000100000; // 1056 0.2577010989189148
storage[794] = -13'b0000100001101; // -269 -0.0656425952911377
storage[795] = -13'b0000111101110; // -494 -0.12057255953550339
storage[796] =  13'b0010010011111; // 1183 0.2887430191040039
storage[797] = -13'b0001001010000; // -592 -0.1445353478193283
storage[798] = -13'b0000010011101; // -157 -0.03837687149643898
storage[799] =  13'b0010100100100; // 1316 0.3212890326976776
storage[800] = -13'b0000110101100; // -428 -0.10458045452833176
storage[801] = -13'b0011001111011; // -1659 -0.4049086272716522
storage[802] = -13'b0000001110011; // -115 -0.028102684766054153
storage[803] = -13'b0000010010011; // -147 -0.035917915403842926
storage[804] =  13'b0011011101111; // 1775 0.4332297742366791
storage[805] = -13'b0001001001110; // -590 -0.14399710297584534
storage[806] =  13'b0000001110000; // 112 0.027436355128884315
storage[807] =  13'b0010001011110; // 1118 0.2729060649871826
storage[808] = -13'b0000111111111; // -511 -0.12480736523866653
storage[809] = -13'b0010001000011; // -1091 -0.26645952463150024
storage[810] = -13'b0001011010100; // -724 -0.1768464595079422
storage[811] = -13'b0010001000010; // -1090 -0.266152024269104
storage[812] = -13'b0000101110010; // -370 -0.09039510786533356
storage[813] = -13'b0000000101001; // -41 -0.009979883208870888
storage[814] = -13'b0001000110010; // -562 -0.13723137974739075
storage[815] = -13'b0000001110111; // -119 -0.029140405356884003
storage[816] =  13'b0001100001010; // 778 0.1898335963487625
storage[817] = -13'b0000101011110; // -350 -0.08546406030654907
storage[818] = -13'b0000110010011; // -403 -0.09836436063051224
storage[819] =  13'b0011110101110; // 1966 0.47986090183258057
storage[820] =  13'b0000110101110; // 430 0.10500121116638184
storage[821] =  13'b0001101111011; // 891 0.2175908237695694
storage[822] =  13'b0001111010000; // 976 0.23829324543476105
storage[823] =  13'b0001000011101; // 541 0.1321912556886673
storage[824] =  13'b0001011111000; // 760 0.18548265099525452
storage[825] =  13'b0010000101000; // 1064 0.25971323251724243
storage[826] =  13'b0000100110110; // 310 0.07564359158277512
storage[827] =  13'b0001111011001; // 985 0.24040661752223969
storage[828] =  13'b0001010100010; // 674 0.1645474135875702
storage[829] =  13'b0000001111110; // 126 0.0308048278093338
storage[830] =  13'b0000001001011; // 75 0.01821848936378956
storage[831] = -13'b0000111100001; // -481 -0.11748833954334259
storage[832] =  13'b0000100100000; // 288 0.07028702646493912
storage[833] = -13'b0001001000110; // -582 -0.1421038806438446
storage[834] = -13'b0000101011011; // -347 -0.08478744328022003
storage[835] = -13'b0001010101100; // -684 -0.1670403629541397
storage[836] = -13'b0000110111100; // -444 -0.10846761614084244
storage[837] = -13'b0000110011001; // -409 -0.09996910393238068
storage[838] = -13'b0000100101101; // -301 -0.07359477132558823
storage[839] = -13'b0001110111101; // -957 -0.2335698902606964
storage[840] =  13'b0000011011001; // 217 0.05306718498468399
storage[841] =  13'b0000011010010; // 210 0.051369864493608475
storage[842] = -13'b0001101100100; // -868 -0.21203453838825226
storage[843] = -13'b0000110011111; // -415 -0.10133271664381027
storage[844] =  13'b0000000001110; // 14 0.0033575708512216806
storage[845] = -13'b0000001010010; // -82 -0.019926011562347412
storage[846] = -13'b0000011000110; // -198 -0.04842698201537132
storage[847] = -13'b0000111100001; // -481 -0.11753319203853607
storage[848] = -13'b0010101000101; // -1349 -0.32940468192100525
storage[849] = -13'b0010101110111; // -1399 -0.34150153398513794
storage[850] =  13'b0000010111100; // 188 0.045951005071401596
storage[851] =  13'b0000000100000; // 32 0.007795979268848896
storage[852] =  13'b0000011011101; // 221 0.05401099473237991
storage[853] =  13'b0010001100001; // 1121 0.27359312772750854
storage[854] =  13'b0001101110001; // 881 0.21501855552196503
storage[855] =  13'b0001001100101; // 613 0.14956137537956238
storage[856] =  13'b0000001100011; // 99 0.02410346083343029
storage[857] =  13'b0000000010111; // 23 0.00558395916596055
storage[858] = -13'b0000010011110; // -158 -0.03859752044081688
storage[859] =  13'b0000011110011; // 243 0.05930030345916748
storage[860] =  13'b0000001001110; // 78 0.018928229808807373
storage[861] =  13'b0000011110000; // 240 0.058603499084711075
storage[862] = -13'b0000001110001; // -113 -0.027500808238983154
storage[863] =  13'b0010000110011; // 1075 0.26256778836250305
storage[864] =  13'b0000101001000; // 328 0.08004488050937653
storage[865] =  13'b0000101100011; // 355 0.08670764416456223
storage[866] =  13'b0000010010011; // 147 0.03600895032286644
storage[867] =  13'b0001011101011; // 747 0.18248093128204346
storage[868] =  13'b0001010000011; // 643 0.1568831354379654
storage[869] =  13'b0001000011111; // 543 0.1325596123933792
storage[870] =  13'b0001111111010; // 1018 0.24850480258464813
storage[871] =  13'b0000010101001; // 169 0.04127585515379906
storage[872] =  13'b0001000110110; // 566 0.13811813294887543
storage[873] =  13'b0000101100011; // 355 0.08675592392683029
storage[874] = -13'b0000010011111; // -159 -0.038862451910972595
storage[875] =  13'b0000001111001; // 121 0.029618898406624794
storage[876] = -13'b0001000110001; // -561 -0.13706302642822266
storage[877] = -13'b0000101100111; // -359 -0.08766677975654602
storage[878] = -13'b0010001000001; // -1089 -0.2658117413520813
storage[879] = -13'b0010000110101; // -1077 -0.2630454897880554
storage[880] =  13'b0000100100110; // 294 0.07174696028232574
storage[881] = -13'b0010001001011; // -1099 -0.26826632022857666
storage[882] = -13'b0000110001010; // -394 -0.09612362086772919
storage[883] =  13'b0010010010011; // 1171 0.28588828444480896
storage[884] = -13'b0001000010010; // -530 -0.1294568032026291
storage[885] =  13'b0000101001101; // 333 0.08128770440816879
storage[886] = -13'b0001011110011; // -755 -0.1842537522315979
storage[887] = -13'b0001001000110; // -582 -0.14215052127838135
storage[888] = -13'b0000011111111; // -255 -0.062367234379053116
storage[889] = -13'b0001010110100; // -692 -0.16903546452522278
storage[890] = -13'b0000011110101; // -245 -0.05992323160171509
storage[891] =  13'b0001011101011; // 747 0.18242065608501434
storage[892] = -13'b0001000000101; // -517 -0.12616078555583954
storage[893] = -13'b0000010010111; // -151 -0.03680980205535889
storage[894] =  13'b0001000100001; // 545 0.13295434415340424
storage[895] = -13'b0001101111010; // -890 -0.21737530827522278
storage[896] = -13'b0000011011010; // -218 -0.05331476032733917
storage[897] =  13'b0000000110100; // 52 0.012714946642518044
storage[898] = -13'b0010100001110; // -1294 -0.3159252107143402
storage[899] = -13'b0100001001001; // -2121 -0.517764687538147
storage[900] = -13'b0000100011110; // -286 -0.06993464380502701
storage[901] =  13'b0000001010010; // 82 0.01994241587817669
storage[902] = -13'b0001000011100; // -540 -0.13178622722625732
storage[903] = -13'b0001101111101; // -893 -0.21794280409812927
storage[904] =  13'b0001100011101; // 797 0.19457073509693146
storage[905] = -13'b0000000110000; // -48 -0.011831081472337246
storage[906] =  13'b0000010101001; // 169 0.04121021926403046
storage[907] =  13'b0001110011111; // 927 0.22635330259799957
storage[908] = -13'b0000000110011; // -51 -0.012442616745829582
storage[909] =  13'b0000001011001; // 89 0.02163376286625862
storage[910] = -13'b0001001111010; // -634 -0.15476830303668976
storage[911] =  13'b0000100111111; // 319 0.07792995125055313
storage[912] =  13'b0001000111010; // 570 0.13913662731647491
storage[913] = -13'b0001110000101; // -901 -0.2199457585811615
storage[914] =  13'b0010010001110; // 1166 0.28474995493888855
storage[915] =  13'b0011000011110; // 1566 0.3823060095310211
storage[916] =  13'b0000111111000; // 504 0.12308111041784286
storage[917] =  13'b0010101001111; // 1359 0.3318447768688202
storage[918] =  13'b0001011010001; // 721 0.17600716650485992
storage[919] = -13'b0000011111100; // -252 -0.06150614842772484
storage[920] =  13'b0000111011100; // 476 0.11614184826612473
storage[921] =  13'b0001100001001; // 777 0.18974612653255463
storage[922] =  13'b0010101001010; // 1354 0.33051925897598267
storage[923] =  13'b0000011101101; // 237 0.05794515088200569
storage[924] = -13'b0001000000100; // -516 -0.12606433033943176
storage[925] =  13'b0010100010100; // 1300 0.3173149824142456
storage[926] =  13'b0000010011001; // 153 0.037448134273290634
storage[927] = -13'b0000111101110; // -494 -0.12071500718593597
storage[928] = -13'b0001101000010; // -834 -0.2036186009645462
storage[929] =  13'b0000011101001; // 233 0.056896377354860306
storage[930] =  13'b0000011101011; // 235 0.05741924047470093
storage[931] = -13'b0001001001000; // -584 -0.1426146924495697
storage[932] = -13'b0001010000110; // -646 -0.15778928995132446
storage[933] =  13'b0001101101000; // 872 0.21284307539463043
storage[934] = -13'b0001011001001; // -713 -0.17418871819972992
storage[935] =  13'b0001001100010; // 610 0.14888641238212585
storage[936] =  13'b0000101000110; // 326 0.07970701158046722
storage[937] =  13'b0001010011101; // 669 0.16342902183532715
storage[938] =  13'b0000011110001; // 241 0.05884106084704399
storage[939] = -13'b0000001111010; // -122 -0.02974199317395687
storage[940] = -13'b0000111010011; // -467 -0.11406084895133972
storage[941] =  13'b0000100111010; // 314 0.07677905261516571
storage[942] = -13'b0000111001001; // -457 -0.11154625564813614
storage[943] = -13'b0000110011110; // -414 -0.10096443444490433
storage[944] = -13'b0011101111001; // -1913 -0.4670089781284332
storage[945] =  13'b0000101110101; // 373 0.09105782210826874
storage[946] = -13'b0000000000100; // -4 -0.0009695512126199901
storage[947] = -13'b0000001101000; // -104 -0.02538364566862583
storage[948] = -13'b0001001110111; // -631 -0.15402661263942719
storage[949] = -13'b0001000000111; // -519 -0.12675106525421143
storage[950] = -13'b0000000100000; // -32 -0.00784393586218357
storage[951] =  13'b0000000000010; // 2 0.0003854167298413813
storage[952] = -13'b0000010111111; // -191 -0.046604886651039124
storage[953] = -13'b0101011101101; // -2797 -0.6827574372291565
storage[954] = -13'b0000011010111; // -215 -0.05241220071911812
storage[955] =  13'b0000111001101; // 461 0.11261171847581863
storage[956] =  13'b0000010101011; // 171 0.04183631017804146
storage[957] =  13'b0000001101101; // 109 0.02671814151108265
storage[958] =  13'b0000001101000; // 104 0.025336313992738724
storage[959] =  13'b0000001000110; // 70 0.016990497708320618
storage[960] =  13'b0010001000001; // 1089 0.26589223742485046
storage[961] = -13'b0000110010110; // -406 -0.09909652173519135
storage[962] = -13'b0001100110101; // -821 -0.20044678449630737
storage[963] = -13'b0001010000011; // -643 -0.15694588422775269
storage[964] = -13'b0000101110110; // -374 -0.09137855470180511
storage[965] = -13'b0000110111111; // -447 -0.10905041545629501
storage[966] = -13'b0001100011110; // -798 -0.19487035274505615
storage[967] =  13'b0000110100110; // 422 0.1029813140630722
storage[968] =  13'b0000001110000; // 112 0.027297798544168472
storage[969] = -13'b0010110001010; // -1418 -0.3462189733982086
storage[970] =  13'b0000011100101; // 229 0.0558217391371727
storage[971] =  13'b0000111100110; // 486 0.11863604933023453
storage[972] =  13'b0000000111000; // 56 0.013751933351159096
storage[973] = -13'b0010001100000; // -1120 -0.2734783887863159
storage[974] =  13'b0000010001010; // 138 0.03372731804847717
storage[975] =  13'b0000110010000; // 400 0.097666434943676
storage[976] = -13'b0000010101001; // -169 -0.041158344596624374
storage[977] = -13'b0000110000000; // -384 -0.09363864362239838
storage[978] = -13'b0001101111101; // -893 -0.21798932552337646
storage[979] =  13'b0001011101000; // 744 0.18154990673065186
storage[980] =  13'b0001001101011; // 619 0.15117928385734558
storage[981] = -13'b0001000101101; // -557 -0.13590848445892334
storage[982] = -13'b0000111101000; // -488 -0.1192518025636673
storage[983] = -13'b0000011011100; // -220 -0.053828682750463486
storage[984] = -13'b0011101010101; // -1877 -0.4581741690635681
storage[985] =  13'b0000011011111; // 223 0.05448430776596069
storage[986] =  13'b0000111000110; // 454 0.11075695604085922
storage[987] = -13'b0001000110110; // -566 -0.13823820650577545
storage[988] =  13'b0000101100011; // 355 0.08676862716674805
storage[989] =  13'b0010011011111; // 1247 0.3043883740901947
storage[990] =  13'b0000101110111; // 375 0.09155373275279999
storage[991] =  13'b0000110111000; // 440 0.10742546617984772
storage[992] =  13'b0010110001111; // 1423 0.34730517864227295
storage[993] =  13'b0011011111111; // 1791 0.4373694956302643
storage[994] =  13'b0001111101011; // 1003 0.24487878382205963
storage[995] =  13'b0010010000111; // 1159 0.28299519419670105
storage[996] =  13'b0010001101100; // 1132 0.2762811481952667
storage[997] =  13'b0000011110100; // 244 0.059476010501384735
storage[998] =  13'b0000011011110; // 222 0.05428321287035942
storage[999] = -13'b0011010111011; // -1723 -0.42070960998535156
storage[1000] = -13'b0000001011110; // -94 -0.022923899814486504
storage[1001] = -13'b0000101100101; // -357 -0.08724183589220047
storage[1002] = -13'b0001101010001; // -849 -0.20716553926467896
storage[1003] =  13'b0001001001001; // 585 0.1427905112504959
storage[1004] = -13'b0001101011000; // -856 -0.20889493823051453
storage[1005] = -13'b0010001010101; // -1109 -0.2708547115325928
storage[1006] =  13'b0000101111110; // 382 0.0933210626244545
storage[1007] = -13'b0000101101110; // -366 -0.08934587985277176
storage[1008] = -13'b0010100110001; // -1329 -0.32455745339393616
storage[1009] =  13'b0000011000010; // 194 0.047298282384872437
storage[1010] = -13'b0000000010111; // -23 -0.005562592763453722
storage[1011] =  13'b0001000000001; // 513 0.12531881034374237
storage[1012] =  13'b0000001111111; // 127 0.03105301968753338
storage[1013] = -13'b0000110110100; // -436 -0.1065104529261589
storage[1014] =  13'b0000110010100; // 404 0.09854330122470856
storage[1015] =  13'b0001000011111; // 543 0.13263048231601715
storage[1016] = -13'b0001010011000; // -664 -0.16209575533866882
storage[1017] = -13'b0000110010110; // -406 -0.0991533100605011
storage[1018] = -13'b0000011010101; // -213 -0.051887694746255875
storage[1019] =  13'b0000011000111; // 199 0.04855829477310181
storage[1020] =  13'b0000001100110; // 102 0.024971481412649155
storage[1021] =  13'b0010011101111; // 1263 0.30838289856910706
storage[1022] =  13'b0000000010110; // 22 0.005444343667477369
storage[1023] =  13'b0000001111100; // 124 0.030154692009091377
storage[1024] =  13'b0000111001011; // 459 0.11199090629816055
storage[1025] = -13'b0000110010011; // -403 -0.09850437194108963
storage[1026] = -13'b0001110100011; // -931 -0.2272663116455078
storage[1027] =  13'b0001101011101; // 861 0.21032153069972992
storage[1028] =  13'b0001000101000; // 552 0.13487474620342255
storage[1029] =  13'b0011000000010; // 1538 0.3754759132862091
storage[1030] =  13'b0001101100011; // 867 0.21167388558387756
storage[1031] =  13'b0010000011011; // 1051 0.2565910220146179
storage[1032] =  13'b0000101000011; // 323 0.07879917323589325
storage[1033] =  13'b0011000010101; // 1557 0.3800594210624695
storage[1034] =  13'b0000001111011; // 123 0.030108533799648285
storage[1035] =  13'b0001011000000; // 704 0.17184709012508392
storage[1036] =  13'b0000010011100; // 156 0.03812061622738838
storage[1037] = -13'b0010000000000; // -1024 -0.24998891353607178
storage[1038] = -13'b0011001011000; // -1624 -0.3965962529182434
storage[1039] = -13'b0000011111111; // -255 -0.06218301132321358
storage[1040] = -13'b0010000100110; // -1062 -0.2592116594314575
storage[1041] =  13'b0000000101101; // 45 0.011098109185695648
storage[1042] = -13'b0000000101001; // -41 -0.01002782303839922
storage[1043] = -13'b0000000000010; // -2 -0.00045431542093865573
storage[1044] = -13'b0000000110010; // -50 -0.012198176234960556
storage[1045] = -13'b0000101000000; // -320 -0.0782390832901001
storage[1046] = -13'b0000010111010; // -186 -0.04539155215024948
storage[1047] =  13'b0001110001111; // 911 0.2225223034620285
storage[1048] =  13'b0000110111011; // 443 0.10814701020717621
storage[1049] =  13'b0010001001110; // 1102 0.2691068649291992
storage[1050] =  13'b0011010011010; // 1690 0.4126179814338684
storage[1051] =  13'b0000110000110; // 390 0.09529032558202744
storage[1052] =  13'b0001101100010; // 866 0.21148069202899933
storage[1053] = -13'b0000010100000; // -160 -0.0389481820166111
storage[1054] =  13'b0000110000011; // 387 0.09454236924648285
storage[1055] = -13'b0001000001110; // -526 -0.1285206526517868
storage[1056] = -13'b0000001011011; // -91 -0.022188562899827957
storage[1057] =  13'b0000111111100; // 508 0.12413787841796875
storage[1058] =  13'b0000101001100; // 332 0.08106997609138489
storage[1059] =  13'b0001000010011; // 531 0.1296631544828415
storage[1060] =  13'b0000100011010; // 282 0.06892979890108109
storage[1061] = -13'b0001000111001; // -569 -0.13902999460697174
storage[1062] = -13'b0000111001011; // -459 -0.11199592053890228
storage[1063] =  13'b0001101000010; // 834 0.2035442739725113
storage[1064] =  13'b0000110111010; // 442 0.10779489576816559
storage[1065] = -13'b0010001100000; // -1120 -0.27348941564559937
storage[1066] = -13'b0000110010011; // -403 -0.09838392585515976
storage[1067] = -13'b0001101100100; // -868 -0.211976557970047
storage[1068] = -13'b0100101111100; // -2428 -0.5926762223243713
storage[1069] = -13'b0000000110001; // -49 -0.012063352391123772
storage[1070] = -13'b0000010100101; // -165 -0.04028952866792679
storage[1071] = -13'b0100001010011; // -2131 -0.5203232765197754
storage[1072] = -13'b0001001101000; // -616 -0.15035131573677063
storage[1073] =  13'b0000111000100; // 452 0.11025969684123993
storage[1074] =  13'b0010010010001; // 1169 0.2854366898536682
storage[1075] =  13'b0000111011111; // 479 0.11693982779979706
storage[1076] =  13'b0000000101110; // 46 0.011271845549345016
storage[1077] =  13'b0000011101101; // 237 0.057950060814619064
storage[1078] =  13'b0000001100010; // 98 0.023886332288384438
storage[1079] = -13'b0000011010010; // -210 -0.0512315072119236
storage[1080] = -13'b0000111110101; // -501 -0.12220890074968338
storage[1081] = -13'b0001011001101; // -717 -0.17500744760036469
storage[1082] = -13'b0011011011101; // -1757 -0.4289860725402832
storage[1083] = -13'b0000100101101; // -301 -0.07355906814336777
storage[1084] = -13'b0010000100111; // -1063 -0.2594415545463562
storage[1085] = -13'b0011010110111; // -1719 -0.419689804315567
storage[1086] = -13'b0001011111100; // -764 -0.18646179139614105
storage[1087] =  13'b0001100001000; // 776 0.18950024247169495
storage[1088] =  13'b0010000000100; // 1028 0.2509863078594208
storage[1089] =  13'b0000010011001; // 153 0.03743183985352516
storage[1090] =  13'b0001101011101; // 861 0.2101842314004898
storage[1091] =  13'b0000111010101; // 469 0.11452911794185638
storage[1092] =  13'b0001010110111; // 695 0.1696900874376297
storage[1093] = -13'b0000000011000; // -24 -0.005744146183133125
storage[1094] =  13'b0000110100111; // 423 0.10329542309045792
storage[1095] =  13'b0001001001010; // 586 0.14308181405067444
storage[1096] =  13'b0000010100011; // 163 0.03984362259507179
storage[1097] = -13'b0001011100101; // -741 -0.1808525174856186
storage[1098] =  13'b0000110100011; // 419 0.10231926292181015
storage[1099] = -13'b0000010010110; // -150 -0.03660022094845772
storage[1100] =  13'b0001100011000; // 792 0.1934613585472107
storage[1101] = -13'b0000101111001; // -377 -0.09205587208271027
storage[1102] =  13'b0010011010111; // 1239 0.30250856280326843
storage[1103] =  13'b0001111110001; // 1009 0.2462867647409439
storage[1104] = -13'b0000000001001; // -9 -0.0022181831300258636
storage[1105] =  13'b0010010001010; // 1162 0.28362780809402466
storage[1106] = -13'b0000100000010; // -258 -0.06296173483133316
storage[1107] =  13'b0000010101111; // 175 0.04281022772192955
storage[1108] =  13'b0001100010100; // 788 0.19241322576999664
storage[1109] = -13'b0000000110011; // -51 -0.012545476667582989
storage[1110] =  13'b0001011011101; // 733 0.17892736196517944
storage[1111] =  13'b0010011000110; // 1222 0.2984389066696167
storage[1112] = -13'b0001101101000; // -872 -0.2129768431186676
storage[1113] = -13'b0001110001000; // -904 -0.22061218321323395
storage[1114] =  13'b0010000000010; // 1026 0.2503851056098938
storage[1115] = -13'b0010010011110; // -1182 -0.288628488779068
storage[1116] = -13'b0001111011111; // -991 -0.24202822148799896
storage[1117] = -13'b0001000111111; // -575 -0.14033755660057068
storage[1118] =  13'b0000010110001; // 177 0.04321199283003807
storage[1119] =  13'b0000000001010; // 10 0.002401186851784587
storage[1120] =  13'b0000010000111; // 135 0.032840944826602936
storage[1121] =  13'b0001001100110; // 614 0.14978565275669098
storage[1122] =  13'b0000001100111; // 103 0.025052599608898163
storage[1123] =  13'b0001001110101; // 629 0.15347376465797424
storage[1124] =  13'b0001110111000; // 952 0.232540562748909
storage[1125] =  13'b0001110011100; // 924 0.22557906806468964
storage[1126] =  13'b0001101101101; // 877 0.21418003737926483
storage[1127] =  13'b0001011110010; // 754 0.1841648668050766
storage[1128] =  13'b0001011110110; // 758 0.18502095341682434
storage[1129] = -13'b0001110111000; // -952 -0.23245786130428314
storage[1130] =  13'b0000011011010; // 218 0.05318703502416611
storage[1131] =  13'b0001001011011; // 603 0.14732012152671814
storage[1132] = -13'b0010011111101; // -1277 -0.3116615116596222
storage[1133] = -13'b0001010100011; // -675 -0.164829820394516
storage[1134] =  13'b0000001011100; // 92 0.022565091028809547
storage[1135] = -13'b0010010110111; // -1207 -0.2946023643016815
storage[1136] = -13'b0101001111100; // -2684 -0.6553308963775635
storage[1137] = -13'b0101001000011; // -2627 -0.6413962841033936
storage[1138] = -13'b0000010010100; // -148 -0.03607990965247154
storage[1139] = -13'b0011011111000; // -1784 -0.4355463981628418
storage[1140] = -13'b0011011011100; // -1756 -0.4287988245487213
storage[1141] =  13'b0001011001011; // 715 0.17468218505382538
storage[1142] = -13'b0011100101100; // -1836 -0.4482119679450989
storage[1143] = -13'b0001110000101; // -901 -0.2198835015296936
storage[1144] =  13'b0000101110100; // 372 0.09091944992542267
storage[1145] =  13'b0000010101110; // 174 0.04246026277542114
storage[1146] = -13'b0000101000000; // -320 -0.07804340869188309
storage[1147] =  13'b0000010010111; // 151 0.03679913654923439
storage[1148] =  13'b0001000101111; // 559 0.13638712465763092
storage[1149] = -13'b0000101111001; // -377 -0.09205193817615509
storage[1150] = -13'b0000010111100; // -188 -0.04580763354897499
storage[1151] =  13'b0001000111010; // 570 0.13917818665504456
storage[1152] =  13'b0010101100011; // 1379 0.33660688996315
storage[1153] =  13'b0001010001001; // 649 0.15840782225131989
storage[1154] = -13'b0000101001011; // -331 -0.0807914212346077
storage[1155] = -13'b0000010110011; // -179 -0.043705400079488754
storage[1156] =  13'b0001111100100; // 996 0.243256613612175
storage[1157] = -13'b0001000001010; // -522 -0.12740127742290497
storage[1158] = -13'b0000001010000; // -80 -0.019483497366309166
storage[1159] = -13'b0010100101010; // -1322 -0.322681188583374
storage[1160] = -13'b0000011101011; // -235 -0.05727381259202957
storage[1161] = -13'b0000000000111; // -7 -0.0016551731387153268
storage[1162] =  13'b0001100001001; // 777 0.18963010609149933
storage[1163] =  13'b0000011010110; // 214 0.05222995579242706
storage[1164] =  13'b0000110000101; // 389 0.0949300080537796
storage[1165] =  13'b0000000010011; // 19 0.004677562974393368
storage[1166] =  13'b0000001000101; // 69 0.016873685643076897
storage[1167] = -13'b0000011011100; // -220 -0.05371639505028725
storage[1168] = -13'b0000011010101; // -213 -0.05200354754924774
storage[1169] =  13'b0000010010010; // 146 0.03570708632469177
storage[1170] = -13'b0001001011101; // -605 -0.14773514866828918
storage[1171] = -13'b0001001110011; // -627 -0.15300939977169037
storage[1172] = -13'b0001100010000; // -784 -0.1913248896598816
storage[1173] = -13'b0000110001000; // -392 -0.09569652378559113
storage[1174] = -13'b0010101101011; // -1387 -0.3387351334095001
storage[1175] = -13'b0011000010101; // -1557 -0.38019993901252747
storage[1176] = -13'b0010100100000; // -1312 -0.3203445076942444
storage[1177] = -13'b0000101100001; // -353 -0.08609703183174133
storage[1178] = -13'b0000001100000; // -96 -0.023417510092258453
storage[1179] = -13'b0000000000111; // -7 -0.0017526772571727633
storage[1180] = -13'b0010001010101; // -1109 -0.27086135745048523
storage[1181] = -13'b0001001110100; // -628 -0.15329591929912567
storage[1182] =  13'b0001011111000; // 760 0.18565557897090912
storage[1183] = -13'b0000001101100; // -108 -0.026373783126473427
storage[1184] = -13'b0001001000010; // -578 -0.14100609719753265
storage[1185] =  13'b0001000001011; // 523 0.12777887284755707
storage[1186] = -13'b0000111100010; // -482 -0.11756712943315506
storage[1187] = -13'b0010101000110; // -1350 -0.3296218514442444
storage[1188] =  13'b0001000100000; // 544 0.132846400141716
storage[1189] =  13'b0000001111000; // 120 0.029369529336690903
storage[1190] =  13'b0001000100100; // 548 0.13383522629737854
storage[1191] = -13'b0000110010000; // -400 -0.09762464463710785
storage[1192] = -13'b0000101010000; // -336 -0.08202461898326874
storage[1193] = -13'b0000000100101; // -37 -0.009133563376963139
storage[1194] = -13'b0000011110001; // -241 -0.05886033922433853
storage[1195] =  13'b0010100100001; // 1313 0.3206437826156616
storage[1196] = -13'b0000011100011; // -227 -0.055427998304367065
storage[1197] = -13'b0000100101111; // -303 -0.07402042299509048
storage[1198] = -13'b0000011111001; // -249 -0.060827672481536865
storage[1199] =  13'b0000000111101; // 61 0.014964166097342968
storage[1200] =  13'b0000100000100; // 260 0.0634758472442627
storage[1201] = -13'b0000001011101; // -93 -0.022662026807665825
storage[1202] =  13'b0001110101001; // 937 0.22881977260112762
storage[1203] =  13'b0001111001000; // 968 0.236276775598526
storage[1204] =  13'b0000101110101; // 373 0.09114940464496613
storage[1205] =  13'b0010111111111; // 1535 0.37463468313217163
storage[1206] =  13'b0000001101100; // 108 0.02636718563735485
storage[1207] =  13'b0000000111100; // 60 0.014611811377108097
storage[1208] = -13'b0010100100111; // -1319 -0.3220764994621277
storage[1209] = -13'b0000101100000; // -352 -0.08589412271976471
storage[1210] = -13'b0001010101111; // -687 -0.16764923930168152
storage[1211] = -13'b0010011101101; // -1261 -0.30790868401527405
storage[1212] = -13'b0011100010011; // -1811 -0.4421943724155426
storage[1213] =  13'b0001010001001; // 649 0.1585296392440796
storage[1214] = -13'b0001011101000; // -744 -0.1816018968820572
storage[1215] =  13'b0000011101010; // 234 0.057199377566576004
storage[1216] =  13'b0000100011101; // 285 0.06947112828493118
storage[1217] = -13'b0001000010000; // -528 -0.12881268560886383
storage[1218] =  13'b0001111001010; // 970 0.2368449866771698
storage[1219] =  13'b0001010101000; // 680 0.16590861976146698
storage[1220] =  13'b0010000000011; // 1027 0.25061145424842834
storage[1221] =  13'b0010101011100; // 1372 0.3350025713443756
storage[1222] = -13'b0000000011100; // -28 -0.006828243378549814
storage[1223] = -13'b0001110111101; // -957 -0.23370696604251862
storage[1224] = -13'b0000001000101; // -69 -0.016918525099754333
storage[1225] =  13'b0000000110101; // 53 0.01300840824842453
storage[1226] =  13'b0000011011110; // 222 0.05430680140852928
storage[1227] =  13'b0000100111001; // 313 0.07632080465555191
storage[1228] =  13'b0000011001001; // 201 0.04915311932563782
storage[1229] =  13'b0001011000010; // 706 0.1722526252269745
storage[1230] = -13'b0001000110101; // -565 -0.13789987564086914
storage[1231] =  13'b0000110001000; // 392 0.09576296806335449
storage[1232] =  13'b0000100010111; // 279 0.06815735250711441
storage[1233] =  13'b0000000000001; // 1 0.00018701048975344747
storage[1234] =  13'b0001001100101; // 613 0.14958111941814423
storage[1235] = -13'b0000101100011; // -355 -0.08661852777004242
storage[1236] = -13'b0000010100011; // -163 -0.039841484278440475
storage[1237] = -13'b0000101011110; // -350 -0.08543142676353455
storage[1238] = -13'b0000111100010; // -482 -0.11764194816350937
storage[1239] = -13'b0000011110111; // -247 -0.060271456837654114
storage[1240] =  13'b0000001111010; // 122 0.029723986983299255
storage[1241] =  13'b0001010011110; // 670 0.1635950803756714
storage[1242] = -13'b0000101100001; // -353 -0.08614508807659149
storage[1243] = -13'b0010000001101; // -1037 -0.2532047927379608
storage[1244] = -13'b0011111101010; // -2026 -0.4945346415042877
storage[1245] = -13'b0001111001010; // -970 -0.2368714064359665
storage[1246] = -13'b0000110000101; // -389 -0.09494303911924362
storage[1247] = -13'b0010111001001; // -1481 -0.3616845905780792
storage[1248] =  13'b0001011100011; // 739 0.18036311864852905
storage[1249] =  13'b0001101100010; // 866 0.21131113171577454
storage[1250] = -13'b0000110001101; // -397 -0.09698479622602463
storage[1251] = -13'b0001011001011; // -715 -0.1746320128440857
storage[1252] = -13'b0001100010011; // -787 -0.19215907156467438
storage[1253] = -13'b0010111001011; // -1483 -0.3620096445083618
storage[1254] = -13'b0010111010101; // -1493 -0.36460965871810913
storage[1255] = -13'b0000110010111; // -407 -0.09938806295394897
storage[1256] = -13'b0010100001111; // -1295 -0.3162839710712433
storage[1257] = -13'b0000110110101; // -437 -0.10666552186012268
storage[1258] =  13'b0000011001100; // 204 0.04980985075235367
storage[1259] = -13'b0010100101011; // -1323 -0.3229599893093109
storage[1260] =  13'b0000001000000; // 64 0.015655335038900375
storage[1261] =  13'b0000001111000; // 120 0.02934631146490574
storage[1262] = -13'b0000101110101; // -373 -0.0910477414727211
storage[1263] = -13'b0000000100011; // -35 -0.008586309850215912
storage[1264] = -13'b0000101100110; // -358 -0.08731400966644287
storage[1265] = -13'b0000011110011; // -243 -0.05938419699668884
storage[1266] = -13'b0000010000111; // -135 -0.033048857003450394
storage[1267] = -13'b0000010110101; // -181 -0.04410815238952637
storage[1268] =  13'b0001000000101; // 517 0.12629473209381104
storage[1269] = -13'b0000011101011; // -235 -0.057416267693042755
storage[1270] = -13'b0001010111011; // -699 -0.17064866423606873
storage[1271] =  13'b0000001111110; // 126 0.030690476298332214
storage[1272] =  13'b0001000101011; // 555 0.13552431762218475
storage[1273] =  13'b0001000010111; // 535 0.13062018156051636
storage[1274] =  13'b0000110000001; // 385 0.09389291703701019
storage[1275] =  13'b0000110001110; // 398 0.09708062559366226
storage[1276] =  13'b0000111000000; // 448 0.10946966707706451
storage[1277] =  13'b0000110110001; // 433 0.1056002825498581
storage[1278] =  13'b0000111001010; // 458 0.11192923039197922
storage[1279] =  13'b0000101110100; // 372 0.09087169915437698
storage[1280] = -13'b0000010001010; // -138 -0.03369428217411041
storage[1281] = -13'b0010000000111; // -1031 -0.2517126500606537
storage[1282] = -13'b0001010001010; // -650 -0.15879632532596588
storage[1283] = -13'b0001000101011; // -555 -0.13557370007038116
storage[1284] = -13'b0000000111011; // -59 -0.014312735758721828
storage[1285] = -13'b0010100001011; // -1291 -0.31527817249298096
storage[1286] = -13'b0001001110100; // -628 -0.1532008945941925
storage[1287] = -13'b0000010110000; // -176 -0.042999204248189926
storage[1288] = -13'b0000110001001; // -393 -0.09583450108766556
storage[1289] =  13'b0000010111011; // 187 0.0456157885491848
storage[1290] =  13'b0001101011100; // 860 0.21005460619926453
storage[1291] = -13'b0000011010010; // -210 -0.05131220072507858
storage[1292] =  13'b0000010110000; // 176 0.042897410690784454
storage[1293] =  13'b0001000100111; // 551 0.1345868855714798
storage[1294] =  13'b0000000111000; // 56 0.013664772734045982
storage[1295] =  13'b0000100101000; // 296 0.072247713804245
storage[1296] =  13'b0000100000000; // 256 0.062454864382743835
storage[1297] = -13'b0000100010001; // -273 -0.06677154451608658
storage[1298] =  13'b0000000011001; // 25 0.006109831854701042
storage[1299] =  13'b0000100000001; // 257 0.0627775490283966
storage[1300] = -13'b0000000100110; // -38 -0.009313840419054031
storage[1301] = -13'b0000100101111; // -303 -0.07386071234941483
storage[1302] = -13'b0000001110011; // -115 -0.028171150013804436
storage[1303] =  13'b0000001011001; // 89 0.02178966999053955
storage[1304] = -13'b0000000110101; // -53 -0.012919669970870018
storage[1305] =  13'b0000100000000; // 256 0.06245456263422966
storage[1306] = -13'b0001101010000; // -848 -0.20693480968475342
storage[1307] = -13'b0000000111010; // -58 -0.014054100960493088
storage[1308] = -13'b0000010001001; // -137 -0.033460844308137894
storage[1309] = -13'b0000101111110; // -382 -0.09327895939350128
storage[1310] =  13'b0000001001101; // 77 0.01879267767071724
storage[1311] =  13'b0000100101100; // 300 0.07319096475839615
storage[1312] = -13'b0000010111111; // -191 -0.04665647819638252
storage[1313] =  13'b0000100000100; // 260 0.06340982019901276
storage[1314] =  13'b0000111111010; // 506 0.12341571599245071
storage[1315] = -13'b0000010111001; // -185 -0.045122645795345306
storage[1316] = -13'b0000001111101; // -125 -0.030467592179775238
storage[1317] =  13'b0001101010001; // 849 0.20726053416728973
storage[1318] = -13'b0000010011011; // -155 -0.03792506828904152
storage[1319] =  13'b0000000111101; // 61 0.014906959608197212
storage[1320] =  13'b0001000010011; // 531 0.12966148555278778
storage[1321] =  13'b0000101000010; // 322 0.07851456105709076
storage[1322] =  13'b0000010001010; // 138 0.033642783761024475
storage[1323] = -13'b0000000111101; // -61 -0.014972774311900139
storage[1324] = -13'b0001101101001; // -873 -0.21309475600719452
storage[1325] = -13'b0001101001001; // -841 -0.20527327060699463
storage[1326] = -13'b0000001011001; // -89 -0.021668359637260437
storage[1327] = -13'b0010100000100; // -1284 -0.3133620321750641
storage[1328] = -13'b0001101000001; // -833 -0.20333555340766907
storage[1329] = -13'b0000110110110; // -438 -0.106834776699543
storage[1330] = -13'b0011100000010; // -1794 -0.4380530118942261
storage[1331] = -13'b0001011011001; // -729 -0.17793765664100647
storage[1332] =  13'b0001010110110; // 694 0.16935056447982788
storage[1333] = -13'b0100100010011; // -2323 -0.5670378804206848
storage[1334] = -13'b0011000101000; // -1576 -0.38468289375305176
storage[1335] = -13'b0000011000110; // -198 -0.048431482166051865
storage[1336] = -13'b0011110110110; // -1974 -0.4819732904434204
storage[1337] =  13'b0000101010011; // 339 0.08284606039524078
storage[1338] =  13'b0001011110010; // 754 0.18401479721069336
storage[1339] =  13'b0000011000110; // 198 0.04822491854429245
storage[1340] =  13'b0000110111000; // 440 0.10731470584869385
storage[1341] = -13'b0000011101001; // -233 -0.05688358470797539
storage[1342] =  13'b0000011010001; // 209 0.050937797874212265
storage[1343] =  13'b0000011000000; // 192 0.0469321683049202
storage[1344] = -13'b0001111011101; // -989 -0.24151964485645294
storage[1345] =  13'b0000111001111; // 463 0.11306719481945038
storage[1346] = -13'b0000011111110; // -254 -0.06202143058180809
storage[1347] = -13'b0000100101100; // -300 -0.07323042303323746
storage[1348] = -13'b0000010011101; // -157 -0.03839903324842453
storage[1349] = -13'b0001001001000; // -584 -0.142566978931427
storage[1350] =  13'b0000100110101; // 309 0.07550390064716339
storage[1351] =  13'b0000011101110; // 238 0.05819222703576088
storage[1352] =  13'b0000000111000; // 56 0.013722010888159275
storage[1353] = -13'b0000001001011; // -75 -0.018270809203386307
storage[1354] = -13'b0001111000011; // -963 -0.23507243394851685
storage[1355] = -13'b0000000110011; // -51 -0.012521498836576939
storage[1356] =  13'b0000100001010; // 266 0.06486579030752182
storage[1357] = -13'b0000110000011; // -387 -0.09442145377397537
storage[1358] =  13'b0000101001111; // 335 0.08178169280290604
storage[1359] = -13'b0000100010000; // -272 -0.06641903519630432
storage[1360] = -13'b0001001011101; // -605 -0.14759193360805511
storage[1361] =  13'b0000101100010; // 354 0.0863511934876442
storage[1362] =  13'b0000100110010; // 306 0.07464522868394852
storage[1363] = -13'b0000010011101; // -157 -0.038209401071071625
storage[1364] =  13'b0001011101101; // 749 0.18277227878570557
storage[1365] = -13'b0000100110100; // -308 -0.07528580725193024
storage[1366] =  13'b0000001011100; // 92 0.022394347935914993
storage[1367] = -13'b0000001001110; // -78 -0.01913701742887497
storage[1368] = -13'b0001011001110; // -718 -0.1753283441066742
storage[1369] = -13'b0000000101001; // -41 -0.009893743321299553
storage[1370] =  13'b0000000111110; // 62 0.015208682045340538
storage[1371] = -13'b0000100100100; // -292 -0.07129468023777008
storage[1372] =  13'b0000000100001; // 33 0.008175358176231384
storage[1373] =  13'b0000000101000; // 40 0.009767202660441399
storage[1374] =  13'b0000010011100; // 156 0.03808318451046944
storage[1375] =  13'b0001101001000; // 840 0.2051548808813095
storage[1376] =  13'b0000110100011; // 419 0.10224385559558868
storage[1377] =  13'b0000010010010; // 146 0.03561526536941528
storage[1378] = -13'b0001111100011; // -995 -0.24285587668418884
storage[1379] =  13'b0000010101001; // 169 0.041187819093465805
storage[1380] = -13'b0000000010010; // -18 -0.004491872154176235
storage[1381] =  13'b0000000101010; // 42 0.010348491370677948
storage[1382] =  13'b0000110110010; // 434 0.105929434299469
storage[1383] = -13'b0000010100110; // -166 -0.0405769944190979
storage[1384] =  13'b0001110111010; // 954 0.2329777628183365
storage[1385] =  13'b0000011000111; // 199 0.048499226570129395
storage[1386] = -13'b0000111001000; // -456 -0.11125042289495468
storage[1387] = -13'b0000111001010; // -458 -0.11170408129692078
storage[1388] =  13'b0000101100011; // 355 0.08675230294466019
storage[1389] =  13'b0000001100101; // 101 0.02476854808628559
storage[1390] =  13'b0001000101010; // 554 0.13533887267112732
storage[1391] =  13'b0001010110010; // 690 0.16836968064308167
storage[1392] = -13'b0001000100011; // -547 -0.13343124091625214
storage[1393] =  13'b0000101000110; // 326 0.07956922054290771
storage[1394] = -13'b0000111001011; // -459 -0.1121334508061409
storage[1395] = -13'b0010010000001; // -1153 -0.28148114681243896
storage[1396] = -13'b0001000000110; // -518 -0.12647496163845062
storage[1397] = -13'b0000011001111; // -207 -0.05056387931108475
storage[1398] = -13'b0010000101101; // -1069 -0.2609401345252991
storage[1399] = -13'b0000110100001; // -417 -0.10173157602548599
storage[1400] =  13'b0000100101110; // 302 0.07374565303325653
storage[1401] = -13'b0000100110111; // -311 -0.07598844170570374
storage[1402] = -13'b0000010001010; // -138 -0.033785633742809296
storage[1403] =  13'b0001001101111; // 623 0.1520555019378662
storage[1404] = -13'b0000001001101; // -77 -0.018741656094789505
storage[1405] =  13'b0001010000000; // 640 0.15620116889476776
storage[1406] =  13'b0000011011111; // 223 0.05438968539237976
storage[1407] =  13'b0000011100101; // 229 0.055922385305166245
storage[1408] =  13'b0000001010001; // 81 0.01974533498287201
storage[1409] =  13'b0000011101011; // 235 0.05730360001325607
storage[1410] =  13'b0001001010000; // 592 0.14453180134296417
storage[1411] =  13'b0000100001100; // 268 0.06536798179149628
storage[1412] =  13'b0000100100000; // 288 0.07020916789770126
storage[1413] = -13'b0000110100100; // -420 -0.10263347625732422
storage[1414] = -13'b0000011110101; // -245 -0.05986028164625168
storage[1415] = -13'b0000001000001; // -65 -0.015797939151525497
storage[1416] = -13'b0001000100001; // -545 -0.1331436038017273
storage[1417] =  13'b0000111011010; // 474 0.11564330011606216
storage[1418] = -13'b0000001111011; // -123 -0.030000140890479088
storage[1419] = -13'b0000001000000; // -64 -0.015567519702017307
storage[1420] =  13'b0000011000001; // 193 0.04700164869427681
storage[1421] =  13'b0000001110111; // 119 0.028934231027960777
storage[1422] =  13'b0000010011001; // 153 0.03740251064300537
storage[1423] = -13'b0000011000100; // -196 -0.047810181975364685
storage[1424] = -13'b0000001001011; // -75 -0.01831790618598461
storage[1425] =  13'b0000100101011; // 299 0.07305703312158585
storage[1426] = -13'b0000001010100; // -84 -0.020585883408784866
storage[1427] =  13'b0000011011001; // 217 0.05297162011265755
storage[1428] =  13'b0000011011010; // 218 0.0532430000603199
storage[1429] =  13'b0000010011101; // 157 0.038253676146268845
storage[1430] =  13'b0000101000011; // 323 0.07880307734012604
storage[1431] =  13'b0000100101000; // 296 0.07215524464845657
storage[1432] =  13'b0000010111011; // 187 0.04574384540319443
storage[1433] = -13'b0000100011101; // -285 -0.06953226774930954
storage[1434] = -13'b0001011011011; // -731 -0.17856983840465546
storage[1435] =  13'b0000010000101; // 133 0.032446447759866714
storage[1436] =  13'b0000010110110; // 182 0.04438336566090584
storage[1437] = -13'b0001111110000; // -1008 -0.24601593613624573
storage[1438] = -13'b0000000111011; // -59 -0.01443087961524725
storage[1439] = -13'b0000010101101; // -173 -0.04235532134771347
storage[1440] = -13'b0010100000110; // -1286 -0.3140636682510376
storage[1441] =  13'b0000101100011; // 355 0.08665765076875687
storage[1442] =  13'b0000001101001; // 105 0.025629665702581406
storage[1443] = -13'b0000000000111; // -7 -0.0017966292798519135
storage[1444] =  13'b0000101001010; // 330 0.08047729730606079
storage[1445] =  13'b0000100000111; // 263 0.0641307681798935
storage[1446] = -13'b0000110001011; // -395 -0.09653408825397491
storage[1447] =  13'b0001011011010; // 730 0.17825263738632202
storage[1448] =  13'b0000110010001; // 401 0.09796921908855438
storage[1449] = -13'b0000000001010; // -10 -0.002433560322970152
storage[1450] =  13'b0000011111100; // 252 0.061505500227212906
storage[1451] =  13'b0000000000110; // 6 0.0013446396915242076
storage[1452] =  13'b0000000000010; // 2 0.000559707754291594
storage[1453] =  13'b0000111011001; // 473 0.11540687829256058
storage[1454] =  13'b0000100000110; // 262 0.06403016299009323
storage[1455] = -13'b0000101100100; // -356 -0.08694861829280853
storage[1456] =  13'b0001000000101; // 517 0.12619264423847198
storage[1457] =  13'b0000110000010; // 386 0.09432381391525269
storage[1458] = -13'b0000110000110; // -390 -0.09530371427536011
storage[1459] = -13'b0000000011110; // -30 -0.007372892927378416
storage[1460] = -13'b0000011000111; // -199 -0.0485583059489727
storage[1461] = -13'b0000101010100; // -340 -0.08300721645355225
storage[1462] =  13'b0000010110011; // 179 0.043608248233795166
storage[1463] = -13'b0000010001100; // -140 -0.03419237956404686
storage[1464] = -13'b0001111101110; // -1006 -0.2455347627401352
storage[1465] = -13'b0000010010010; // -146 -0.035583123564720154
storage[1466] = -13'b0001010010101; // -661 -0.16125524044036865
storage[1467] =  13'b0000001110100; // 116 0.028217008337378502
storage[1468] = -13'b0000000100101; // -37 -0.009090450592339039
storage[1469] =  13'b0001011010110; // 726 0.17719729244709015
storage[1470] = -13'b0000000111011; // -59 -0.014502127654850483
storage[1471] = -13'b0000100100011; // -291 -0.07103835791349411
storage[1472] =  13'b0001001111111; // 639 0.15597385168075562
storage[1473] = -13'b0000111010000; // -464 -0.11323200911283493
storage[1474] = -13'b0000110101001; // -425 -0.10381533205509186
storage[1475] =  13'b0000001100001; // 97 0.02377135492861271
storage[1476] =  13'b0000010000001; // 129 0.031563084572553635
storage[1477] =  13'b0000110100111; // 423 0.10334289819002151
storage[1478] =  13'b0000001111101; // 125 0.030614405870437622
storage[1479] =  13'b0000110010000; // 400 0.0975925400853157
storage[1480] =  13'b0000100011110; // 286 0.06976994127035141
storage[1481] =  13'b0000010100000; // 160 0.039030104875564575
storage[1482] =  13'b0000110000110; // 390 0.09509646147489548
storage[1483] = -13'b0000100111000; // -312 -0.07613785564899445
storage[1484] = -13'b0001011010101; // -725 -0.1769404262304306
storage[1485] = -13'b0000010111110; // -190 -0.046441663056612015
storage[1486] =  13'b0000110001011; // 395 0.0964113250374794
storage[1487] =  13'b0001001101101; // 621 0.15171362459659576
storage[1488] =  13'b0000011011111; // 223 0.054452624171972275
storage[1489] =  13'b0000100000100; // 260 0.0635487288236618
storage[1490] =  13'b0001001100101; // 613 0.1496959924697876
storage[1491] =  13'b0000110100101; // 421 0.10271921008825302
storage[1492] = -13'b0000110011001; // -409 -0.09989030659198761
storage[1493] = -13'b0000011010011; // -211 -0.051537662744522095
storage[1494] = -13'b0000011001101; // -205 -0.049973513931035995
storage[1495] =  13'b0000111101000; // 488 0.1190408393740654
storage[1496] = -13'b0000100111011; // -315 -0.0769411027431488
storage[1497] =  13'b0000011001101; // 205 0.05016281083226204
storage[1498] =  13'b0000100011010; // 282 0.06882915645837784
storage[1499] = -13'b0000011101000; // -232 -0.056653570383787155
storage[1500] = -13'b0001011001001; // -713 -0.17409367859363556
storage[1501] =  13'b0000011010101; // 213 0.052088841795921326
storage[1502] = -13'b0000100011001; // -281 -0.0686485767364502
storage[1503] = -13'b0001010111001; // -697 -0.17005276679992676
storage[1504] =  13'b0000011101011; // 235 0.05734262987971306
storage[1505] = -13'b0000001101101; // -109 -0.02649209089577198
storage[1506] = -13'b0000011000100; // -196 -0.0478486530482769
storage[1507] = -13'b0000110110001; // -433 -0.10562998801469803
storage[1508] =  13'b0000001110111; // 119 0.028964834287762642
storage[1509] = -13'b0000011111111; // -255 -0.062192581593990326
storage[1510] = -13'b0001111011011; // -987 -0.2409730702638626
storage[1511] = -13'b0001000100110; // -550 -0.13433612883090973
storage[1512] =  13'b0000001110011; // 115 0.02803991176187992
storage[1513] =  13'b0000010011011; // 155 0.037834830582141876
storage[1514] =  13'b0000011011000; // 216 0.05271657556295395
storage[1515] =  13'b0001000101011; // 555 0.1356019228696823
storage[1516] =  13'b0000000101001; // 41 0.009963244199752808
storage[1517] = -13'b0000000111000; // -56 -0.013613351620733738
storage[1518] =  13'b0000010100010; // 162 0.03943140059709549
storage[1519] = -13'b0000010010101; // -149 -0.03649798780679703
storage[1520] = -13'b0000011010111; // -215 -0.05238688364624977
storage[1521] = -13'b0000000110100; // -52 -0.012624991126358509
storage[1522] =  13'b0000111011010; // 474 0.11571669578552246
storage[1523] =  13'b0000100100001; // 289 0.0706784725189209
storage[1524] =  13'b0000100010111; // 279 0.06817649304866791
storage[1525] =  13'b0000110000010; // 386 0.09421809017658234
storage[1526] =  13'b0001001000000; // 576 0.14068488776683807
storage[1527] =  13'b0001100001001; // 777 0.18972553312778473
storage[1528] = -13'b0001000101001; // -553 -0.13499179482460022
storage[1529] = -13'b0000101110101; // -373 -0.0911659225821495
storage[1530] = -13'b0000100001010; // -266 -0.06483285874128342
storage[1531] =  13'b0000010000000; // 128 0.031137589365243912
storage[1532] =  13'b0000001110100; // 116 0.028227301314473152
storage[1533] =  13'b0001000110000; // 560 0.13660956919193268
storage[1534] = -13'b0000111000100; // -452 -0.11030200123786926
storage[1535] = -13'b0001000000110; // -518 -0.12651808559894562
storage[1536] =  13'b0000000000111; // 7 0.0017770060803741217
storage[1537] = -13'b0001011000110; // -710 -0.17322473227977753
storage[1538] = -13'b0000111100001; // -481 -0.11747890710830688
storage[1539] = -13'b0000101000111; // -327 -0.07987483590841293
storage[1540] = -13'b0000111101011; // -491 -0.11998963356018066
storage[1541] = -13'b0000000111010; // -58 -0.014248287305235863
storage[1542] = -13'b0001010100010; // -674 -0.1644904464483261
storage[1543] =  13'b0000100000111; // 263 0.06420671194791794
storage[1544] = -13'b0000110001110; // -398 -0.09716809540987015
storage[1545] =  13'b0000111011000; // 472 0.11532530933618546
storage[1546] = -13'b0001010100100; // -676 -0.1650000959634781
storage[1547] = -13'b0001101011001; // -857 -0.2093149870634079
storage[1548] = -13'b0000110110011; // -435 -0.1061328649520874
storage[1549] = -13'b0000000010010; // -18 -0.004471155349165201
storage[1550] =  13'b0000000010100; // 20 0.004904015455394983
storage[1551] = -13'b0000011110110; // -246 -0.06009582057595253
storage[1552] = -13'b0000010111010; // -186 -0.0453546978533268
storage[1553] = -13'b0001111111010; // -1018 -0.2486196607351303
storage[1554] = -13'b0010101110100; // -1396 -0.3407266438007355
storage[1555] = -13'b0000000011110; // -30 -0.00743508618324995
storage[1556] = -13'b0000111010100; // -468 -0.11434222012758255
storage[1557] = -13'b0000101000011; // -323 -0.07894609123468399
storage[1558] = -13'b0000010001100; // -140 -0.034265268594026566
storage[1559] =  13'b0000001001001; // 73 0.017893962562084198
storage[1560] =  13'b0000100110000; // 304 0.07425149530172348
storage[1561] =  13'b0000111001101; // 461 0.11257372051477432
storage[1562] =  13'b0000010100000; // 160 0.03906945884227753
storage[1563] =  13'b0000010010100; // 148 0.03616466000676155
storage[1564] = -13'b0001101110101; // -885 -0.21611934900283813
storage[1565] = -13'b0001111000011; // -963 -0.23504386842250824
storage[1566] = -13'b0001001100100; // -612 -0.14944690465927124
storage[1567] = -13'b0001000111001; // -569 -0.13889946043491364
storage[1568] = -13'b0001000111101; // -573 -0.13984353840351105
storage[1569] = -13'b0000100000010; // -258 -0.06306872516870499
storage[1570] = -13'b0000001110010; // -114 -0.027726588770747185
storage[1571] =  13'b0000000110000; // 48 0.011663072742521763
storage[1572] =  13'b0000101011011; // 347 0.08467069268226624
storage[1573] =  13'b0001010110111; // 695 0.1697961986064911
storage[1574] =  13'b0001001110000; // 624 0.15233631432056427
storage[1575] =  13'b0001110000111; // 903 0.2204785943031311
storage[1576] =  13'b0000010101011; // 171 0.04186162352561951
storage[1577] =  13'b0000010110110; // 182 0.04455535486340523
storage[1578] =  13'b0000010010100; // 148 0.036110419780015945
storage[1579] =  13'b0000111001001; // 457 0.1115068569779396
storage[1580] =  13'b0000001000010; // 66 0.016054628416895866
storage[1581] =  13'b0000001100001; // 97 0.023756884038448334
storage[1582] = -13'b0000110110100; // -436 -0.10646932572126389
storage[1583] =  13'b0000100111100; // 316 0.07710904628038406
storage[1584] =  13'b0000111001011; // 459 0.11200663447380066
storage[1585] =  13'b0000001010000; // 80 0.019440623000264168
storage[1586] =  13'b0000001000011; // 67 0.016468405723571777
storage[1587] =  13'b0000001111011; // 123 0.029948793351650238
storage[1588] =  13'b0001011101100; // 748 0.18265053629875183
storage[1589] =  13'b0000101110000; // 368 0.0898299515247345
storage[1590] =  13'b0000010101011; // 171 0.04184954985976219
storage[1591] =  13'b0000101000100; // 324 0.07911866158246994
storage[1592] =  13'b0001000001000; // 520 0.1269691288471222
storage[1593] =  13'b0000100110110; // 310 0.0756395161151886
storage[1594] =  13'b0000010001100; // 140 0.03418547287583351
storage[1595] = -13'b0000000100011; // -35 -0.008598214015364647
storage[1596] = -13'b0000001101100; // -108 -0.026408938691020012
storage[1597] =  13'b0000001000111; // 71 0.017338672652840614
storage[1598] = -13'b0000001001010; // -74 -0.017948243767023087
storage[1599] =  13'b0000000101101; // 45 0.01106178481131792
storage[1600] =  13'b0000000000100; // 4 0.0010409471578896046
storage[1601] = -13'b0000110010100; // -404 -0.09864488244056702
storage[1602] = -13'b0000101011001; // -345 -0.0843423455953598
storage[1603] =  13'b0000000000101; // 5 0.0010987420100718737
storage[1604] =  13'b0000011111111; // 255 0.06222313642501831
storage[1605] = -13'b0000100100101; // -293 -0.07149296253919601
storage[1606] =  13'b0000100010100; // 276 0.06742144376039505
storage[1607] =  13'b0000110000111; // 391 0.09551306068897247
storage[1608] =  13'b0000010101111; // 175 0.04273691028356552
storage[1609] =  13'b0001101000110; // 838 0.20450806617736816
storage[1610] =  13'b0001100100100; // 804 0.19626624882221222
storage[1611] =  13'b0000100111111; // 319 0.07792314141988754
storage[1612] =  13'b0001001110111; // 631 0.15395385026931763
storage[1613] =  13'b0001011011010; // 730 0.17832684516906738
storage[1614] =  13'b0001101001111; // 847 0.20690059661865234
storage[1615] =  13'b0000111000000; // 448 0.10934892296791077
storage[1616] =  13'b0000110011100; // 412 0.10068414360284805
storage[1617] =  13'b0001100011000; // 792 0.1934231072664261
storage[1618] = -13'b0000000101000; // -40 -0.009794934652745724
storage[1619] =  13'b0001010110100; // 692 0.16904287040233612
storage[1620] =  13'b0001101101001; // 873 0.21305087208747864
storage[1621] = -13'b0000111101011; // -491 -0.11978089809417725
storage[1622] = -13'b0000010011111; // -159 -0.03871060535311699
storage[1623] = -13'b0000010000111; // -135 -0.032938189804553986
storage[1624] =  13'b0000110000010; // 386 0.09418189525604248
storage[1625] =  13'b0001000000010; // 514 0.12544327974319458
storage[1626] = -13'b0000010110110; // -182 -0.044539593160152435
storage[1627] =  13'b0000011000011; // 195 0.047589268535375595
storage[1628] =  13'b0000011101010; // 234 0.05709308013319969
storage[1629] =  13'b0001010101100; // 684 0.1670551598072052
storage[1630] =  13'b0000011101011; // 235 0.057455215603113174
storage[1631] =  13'b0000000110101; // 53 0.012834076769649982
storage[1632] =  13'b0000010001110; // 142 0.03473035246133804
storage[1633] =  13'b0000100111111; // 319 0.07793121784925461
storage[1634] =  13'b0000010011010; // 154 0.03748840466141701
storage[1635] = -13'b0000010101011; // -171 -0.041652973741292953
storage[1636] =  13'b0000011010111; // 215 0.052603576332330704
storage[1637] =  13'b0000011001100; // 204 0.04971735179424286
storage[1638] =  13'b0000101100100; // 356 0.08684292435646057
storage[1639] = -13'b0001001010001; // -593 -0.14486092329025269
storage[1640] = -13'b0001000000110; // -518 -0.12656527757644653
storage[1641] = -13'b0000001110000; // -112 -0.027317456901073456
storage[1642] = -13'b0000110101100; // -428 -0.10442518442869186
storage[1643] = -13'b0001100001001; // -777 -0.18963739275932312
storage[1644] = -13'b0001001000101; // -581 -0.14188101887702942
storage[1645] =  13'b0000100001001; // 265 0.06473183631896973
storage[1646] =  13'b0000011000001; // 193 0.047080639749765396
storage[1647] = -13'b0000001000111; // -71 -0.017427267506718636
storage[1648] = -13'b0000101011111; // -351 -0.08564875274896622
storage[1649] = -13'b0000111000010; // -450 -0.10990327596664429
storage[1650] = -13'b0000101001010; // -330 -0.08056505024433136
storage[1651] = -13'b0000011010011; // -211 -0.05143757537007332
storage[1652] = -13'b0000010101110; // -174 -0.04237082228064537
storage[1653] =  13'b0000011001110; // 206 0.05019443482160568
storage[1654] =  13'b0000010101000; // 168 0.04102769121527672
storage[1655] =  13'b0000101111011; // 379 0.09250327944755554
storage[1656] =  13'b0000011100010; // 226 0.055152345448732376
storage[1657] = -13'b0001100011000; // -792 -0.19346819818019867
storage[1658] = -13'b0000010011101; // -157 -0.03824599087238312
storage[1659] = -13'b0000001001100; // -76 -0.018470093607902527
storage[1660] = -13'b0000100011101; // -285 -0.0696120634675026
storage[1661] =  13'b0000001101111; // 111 0.027058107778429985
storage[1662] =  13'b0000111000100; // 452 0.11029884219169617
storage[1663] =  13'b0000010000110; // 134 0.0326872244477272
storage[1664] = -13'b0000000110000; // -48 -0.011699064634740353
storage[1665] =  13'b0000001100001; // 97 0.0236581489443779
storage[1666] = -13'b0000010100110; // -166 -0.04055023193359375
storage[1667] = -13'b0000110100011; // -419 -0.10223518311977386
storage[1668] = -13'b0000100110011; // -307 -0.07493261247873306
storage[1669] = -13'b0001000110001; // -561 -0.13706247508525848
storage[1670] = -13'b0000011011111; // -223 -0.05443008244037628
storage[1671] = -13'b0001010011010; // -666 -0.16257357597351074
storage[1672] =  13'b0000010011010; // 154 0.03748175874352455
storage[1673] =  13'b0000000110011; // 51 0.012497792951762676
storage[1674] =  13'b0000100100100; // 292 0.0713331326842308
storage[1675] = -13'b0000001100011; // -99 -0.02425120770931244
storage[1676] = -13'b0000001000110; // -70 -0.01720123365521431
storage[1677] =  13'b0000011001001; // 201 0.049191053956747055
storage[1678] =  13'b0000010011111; // 159 0.038784801959991455
storage[1679] =  13'b0000000010001; // 17 0.004156269133090973
storage[1680] =  13'b0000101111100; // 380 0.0927494466304779
storage[1681] = -13'b0000000001110; // -14 -0.003398546017706394
storage[1682] = -13'b0000001011100; // -92 -0.022523779422044754
storage[1683] =  13'b0000110001111; // 399 0.09743322432041168
storage[1684] = -13'b0010000110001; // -1073 -0.2620354890823364
storage[1685] = -13'b0010100010000; // -1296 -0.3164535164833069
storage[1686] = -13'b0001110001110; // -910 -0.2220863401889801
storage[1687] = -13'b0000111111111; // -511 -0.12470636516809464
storage[1688] = -13'b0001001100101; // -613 -0.14973647892475128
storage[1689] = -13'b0000100000111; // -263 -0.0642724335193634
storage[1690] = -13'b0001011111000; // -760 -0.18556463718414307
storage[1691] = -13'b0010010011101; // -1181 -0.2882717549800873
storage[1692] = -13'b0000011001000; // -200 -0.04879334196448326
storage[1693] =  13'b0000011010010; // 210 0.051381055265665054
storage[1694] =  13'b0000000110011; // 51 0.012490559369325638
storage[1695] = -13'b0001000001001; // -521 -0.12727871537208557
storage[1696] = -13'b0001000011100; // -540 -0.13188941776752472
storage[1697] = -13'b0000010011010; // -154 -0.037535447627305984
storage[1698] =  13'b0000101110111; // 375 0.09143198281526566
storage[1699] =  13'b0000111011001; // 473 0.11536283791065216
storage[1700] =  13'b0000001010001; // 81 0.019700730219483376
storage[1701] = -13'b0001011100011; // -739 -0.18030866980552673
storage[1702] = -13'b0000011001111; // -207 -0.05054471269249916
storage[1703] =  13'b0000000100000; // 32 0.007781801279634237
storage[1704] = -13'b0000010111100; // -188 -0.0459473617374897
storage[1705] = -13'b0000001011001; // -89 -0.021682314574718475
storage[1706] =  13'b0000011010000; // 208 0.05067836865782738
storage[1707] =  13'b0000011010000; // 208 0.050705622881650925
storage[1708] =  13'b0000000000001; // 1 0.0003183711087331176
storage[1709] = -13'b0000011100111; // -231 -0.05638813599944115
storage[1710] = -13'b0000000010111; // -23 -0.005502961575984955
storage[1711] = -13'b0000010110011; // -179 -0.043736666440963745
storage[1712] = -13'b0000110001100; // -396 -0.09667032212018967
storage[1713] = -13'b0000010100100; // -164 -0.04005811735987663
storage[1714] =  13'b0000011110001; // 241 0.0587284155189991
storage[1715] =  13'b0000010010101; // 149 0.03630431741476059
storage[1716] =  13'b0000100100101; // 293 0.07147836685180664
storage[1717] =  13'b0001110110000; // 944 0.23037824034690857
storage[1718] =  13'b0000110101110; // 430 0.10503216087818146
storage[1719] =  13'b0000010100100; // 164 0.04004376754164696
storage[1720] = -13'b0000100101011; // -299 -0.07290377467870712
storage[1721] = -13'b0001011010111; // -727 -0.17746594548225403
storage[1722] =  13'b0000101101100; // 364 0.08897008746862411
storage[1723] = -13'b0000110100000; // -416 -0.10167085379362106
storage[1724] =  13'b0000000100111; // 39 0.009580360725522041
storage[1725] = -13'b0000001000101; // -69 -0.01695280149579048
storage[1726] = -13'b0000101010001; // -337 -0.08216269314289093
storage[1727] = -13'b0000000101011; // -43 -0.010479808785021305
storage[1728] = -13'b0000010010011; // -147 -0.035855866968631744
storage[1729] = -13'b0000010100011; // -163 -0.039808131754398346
storage[1730] = -13'b0000000000100; // -4 -0.0010526402620598674
storage[1731] =  13'b0000001011110; // 94 0.022984525188803673
storage[1732] =  13'b0000011000110; // 198 0.04832582548260689
storage[1733] =  13'b0000010110011; // 179 0.04359696805477142
storage[1734] =  13'b0000101101001; // 361 0.08812469989061356
storage[1735] =  13'b0000100101010; // 298 0.07285748422145844
storage[1736] = -13'b0000001101100; // -108 -0.026253702118992805
storage[1737] = -13'b0000001010011; // -83 -0.020187409594655037
storage[1738] =  13'b0000011100000; // 224 0.05474628880620003
storage[1739] = -13'b0000011111000; // -248 -0.060462575405836105
storage[1740] =  13'b0001000110100; // 564 0.13760963082313538
storage[1741] =  13'b0000011011001; // 217 0.052980732172727585
storage[1742] =  13'b0001010111100; // 700 0.17082440853118896
storage[1743] =  13'b0001101111110; // 894 0.21833938360214233
storage[1744] =  13'b0001010101010; // 682 0.1665666550397873
storage[1745] =  13'b0000101001111; // 335 0.08179174363613129
storage[1746] =  13'b0000010000000; // 128 0.031226035207509995
storage[1747] = -13'b0000011010100; // -212 -0.05167025700211525
storage[1748] =  13'b0000010011000; // 152 0.037010032683610916
storage[1749] =  13'b0001001101110; // 622 0.15184707939624786
storage[1750] = -13'b0000001000000; // -64 -0.01562913879752159
storage[1751] =  13'b0000000010111; // 23 0.005522990133613348
storage[1752] = -13'b0000010100001; // -161 -0.039201103150844574
storage[1753] =  13'b0000000110011; // 51 0.012516777031123638
storage[1754] = -13'b0000000011001; // -25 -0.006091416347771883
storage[1755] = -13'b0000000100010; // -34 -0.008211668580770493
storage[1756] =  13'b0000000011010; // 26 0.00628064526244998
storage[1757] = -13'b0000001000111; // -71 -0.017370937392115593
storage[1758] = -13'b0000101111001; // -377 -0.09197299182415009
storage[1759] = -13'b0000111110010; // -498 -0.12159261852502823
storage[1760] = -13'b0000010100100; // -164 -0.04012516140937805
storage[1761] =  13'b0000011111010; // 250 0.06096837297081947
storage[1762] =  13'b0000000100001; // 33 0.008037947118282318
storage[1763] =  13'b0000011001110; // 206 0.05021414905786514
storage[1764] =  13'b0000010000100; // 132 0.03224180266261101
storage[1765] = -13'b0000110001101; // -397 -0.09687764942646027
storage[1766] = -13'b0001110010111; // -919 -0.22433525323867798
storage[1767] = -13'b0001010100000; // -672 -0.1640165001153946
storage[1768] =  13'b0000000100010; // 34 0.008310195058584213
storage[1769] = -13'b0001011000010; // -706 -0.17226934432983398
storage[1770] = -13'b0010000100010; // -1058 -0.25818976759910583
storage[1771] = -13'b0000000110100; // -52 -0.012666678987443447
storage[1772] = -13'b0000010001000; // -136 -0.03325101360678673
storage[1773] =  13'b0000111110101; // 501 0.12235935032367706
storage[1774] = -13'b0001111101111; // -1007 -0.24579259753227234
storage[1775] = -13'b0000101000110; // -326 -0.07962065935134888
storage[1776] = -13'b0000000101110; // -46 -0.011227280832827091
storage[1777] = -13'b0000001111010; // -122 -0.02974274568259716
storage[1778] = -13'b0000100110110; // -310 -0.07557803392410278
storage[1779] =  13'b0000000000110; // 6 0.0014382185181602836
storage[1780] =  13'b0000010110011; // 179 0.0437772311270237
storage[1781] = -13'b0000001010110; // -86 -0.021085014566779137
storage[1782] =  13'b0000010011001; // 153 0.03746946156024933
storage[1783] =  13'b0001111100100; // 996 0.2432766705751419
storage[1784] =  13'b0000101011000; // 344 0.08406030386686325
storage[1785] = -13'b0000111011000; // -472 -0.11511717736721039
storage[1786] =  13'b0000110100001; // 417 0.10190355032682419
storage[1787] =  13'b0000111001011; // 459 0.11193934828042984
storage[1788] = -13'b0000110110110; // -438 -0.1068786084651947
storage[1789] =  13'b0000101000111; // 327 0.07993917167186737
storage[1790] =  13'b0000101011100; // 348 0.08493257313966751
storage[1791] =  13'b0001001010000; // 592 0.14442914724349976
storage[1792] =  13'b0000100011001; // 281 0.06850965321063995
storage[1793] =  13'b0000111000010; // 450 0.1098678857088089
storage[1794] =  13'b0000010111001; // 185 0.045285165309906006
storage[1795] =  13'b0001011001110; // 718 0.17533212900161743
storage[1796] =  13'b0010111001011; // 1483 0.36215245723724365
storage[1797] =  13'b0010001010101; // 1109 0.2707379460334778
storage[1798] =  13'b0000011110111; // 247 0.06037557125091553
storage[1799] =  13'b0001011101111; // 751 0.1833924651145935
storage[1800] =  13'b0000111111011; // 507 0.1237923800945282
storage[1801] =  13'b0001001111110; // 638 0.15575002133846283
storage[1802] =  13'b0000111000000; // 448 0.10944916307926178
storage[1803] = -13'b0000001000100; // -68 -0.016531087458133698
storage[1804] = -13'b0000000010111; // -23 -0.005680582486093044
storage[1805] = -13'b0000110100101; // -421 -0.10272570699453354
storage[1806] = -13'b0000110010110; // -406 -0.0991632267832756
storage[1807] =  13'b0001011000000; // 704 0.17180824279785156
storage[1808] =  13'b0000100000000; // 256 0.06250903755426407
storage[1809] =  13'b0000001001100; // 76 0.018516065552830696
storage[1810] =  13'b0000101011001; // 345 0.08433675765991211
storage[1811] =  13'b0000111010100; // 468 0.1143035739660263
storage[1812] = -13'b0000000101101; // -45 -0.010896819643676281
storage[1813] =  13'b0000101010100; // 340 0.08291391283273697
storage[1814] =  13'b0000100000111; // 263 0.06419181078672409
storage[1815] =  13'b0000111001011; // 459 0.11196067929267883
storage[1816] =  13'b0000100101000; // 296 0.07217603921890259
storage[1817] =  13'b0000001111110; // 126 0.030776847153902054
storage[1818] = -13'b0000001011110; // -94 -0.02302926406264305
storage[1819] = -13'b0000011101100; // -236 -0.05764465779066086
storage[1820] = -13'b0000011111100; // -252 -0.0615549236536026
storage[1821] = -13'b0000110001011; // -395 -0.09654232859611511
storage[1822] = -13'b0000011101101; // -237 -0.057909045368433
storage[1823] = -13'b0000011010011; // -211 -0.051436591893434525
storage[1824] = -13'b0000011001010; // -202 -0.04922656714916229
storage[1825] =  13'b0000000010100; // 20 0.004967991262674332
storage[1826] =  13'b0000010101001; // 169 0.04123890772461891
storage[1827] = -13'b0000001111001; // -121 -0.02949994057416916
storage[1828] = -13'b0000001111110; // -126 -0.030736271291971207
storage[1829] = -13'b0000011000011; // -195 -0.047666121274232864
storage[1830] =  13'b0000000010001; // 17 0.004165904596447945
storage[1831] = -13'b0000100000101; // -261 -0.06361857801675797
storage[1832] = -13'b0000000000011; // -3 -0.0006116917938925326
storage[1833] = -13'b0000011010001; // -209 -0.051075488328933716
storage[1834] =  13'b0000011011110; // 222 0.0543065071105957
storage[1835] =  13'b0000011010000; // 208 0.05081065744161606
storage[1836] = -13'b0000100111001; // -313 -0.0764790028333664
storage[1837] =  13'b0000010000001; // 129 0.031582269817590714
storage[1838] = -13'b0000100110110; // -310 -0.07572758942842484
storage[1839] = -13'b0000001011111; // -95 -0.023297986015677452
storage[1840] =  13'b0000000010000; // 16 0.0038209501653909683
storage[1841] = -13'b0000111010001; // -465 -0.11357671022415161
storage[1842] = -13'b0001000110100; // -564 -0.1375880390405655
storage[1843] =  13'b0000000011101; // 29 0.007051789201796055
storage[1844] =  13'b0000110001101; // 397 0.09699372947216034
storage[1845] = -13'b0000011011010; // -218 -0.053147830069065094
storage[1846] = -13'b0000010000111; // -135 -0.03306427225470543
storage[1847] =  13'b0001001011000; // 600 0.14643201231956482
storage[1848] =  13'b0000100001111; // 271 0.06611856073141098
storage[1849] = -13'b0000100011011; // -283 -0.06920409202575684
storage[1850] =  13'b0000101110010; // 370 0.09043273329734802
storage[1851] =  13'b0000000110110; // 54 0.01315415371209383
storage[1852] =  13'b0000100010100; // 276 0.06729237735271454
storage[1853] =  13'b0000110100101; // 421 0.10286971926689148
storage[1854] = -13'b0000010001100; // -140 -0.034160904586315155
storage[1855] = -13'b0000010010011; // -147 -0.0359463095664978
storage[1856] = -13'b0000101011001; // -345 -0.08420342952013016
storage[1857] =  13'b0000011011101; // 221 0.05395174399018288
storage[1858] = -13'b0000101100111; // -359 -0.08770860731601715
storage[1859] =  13'b0000011111011; // 251 0.06121392920613289
storage[1860] =  13'b0000010001010; // 138 0.03380364179611206
storage[1861] =  13'b0000001010100; // 84 0.020505055785179138
storage[1862] =  13'b0000100110010; // 306 0.07480232417583466
storage[1863] = -13'b0000001101010; // -106 -0.025910113006830215
storage[1864] =  13'b0000100001100; // 268 0.06534159928560257
storage[1865] = -13'b0000101011000; // -344 -0.08403022587299347
storage[1866] = -13'b0010101010001; // -1361 -0.3322642147541046
storage[1867] =  13'b0000001110001; // 113 0.027652021497488022
storage[1868] = -13'b0001100110110; // -822 -0.2007303386926651
storage[1869] = -13'b0010110110000; // -1456 -0.3555801212787628
storage[1870] =  13'b0001000011001; // 537 0.13116984069347382
storage[1871] = -13'b0000111010100; // -468 -0.11434558779001236
storage[1872] = -13'b0001001000010; // -578 -0.14107288420200348
storage[1873] =  13'b0000100010001; // 273 0.06666570156812668
storage[1874] = -13'b0000001011101; // -93 -0.022645313292741776
storage[1875] = -13'b0000000111010; // -58 -0.014059040695428848
storage[1876] =  13'b0000101100011; // 355 0.08659495413303375
storage[1877] =  13'b0001000110001; // 561 0.1370353400707245
storage[1878] = -13'b0000001000110; // -70 -0.01720859296619892
storage[1879] =  13'b0000110111111; // 447 0.10921061784029007
storage[1880] =  13'b0000111010111; // 471 0.11499379575252533
storage[1881] = -13'b0000000000111; // -7 -0.0016786260530352592
storage[1882] = -13'b0000001000101; // -69 -0.016953885555267334
storage[1883] = -13'b0000000100100; // -36 -0.00879628211259842
storage[1884] = -13'b0000010010001; // -145 -0.035500623285770416
storage[1885] = -13'b0000001011111; // -95 -0.02328530326485634
storage[1886] = -13'b0000100010001; // -273 -0.06673195213079453
storage[1887] =  13'b0000001100000; // 96 0.023348215967416763
storage[1888] =  13'b0000101100110; // 358 0.08750477433204651
storage[1889] =  13'b0000010101111; // 175 0.04278135299682617
storage[1890] =  13'b0000010111011; // 187 0.045570164918899536
storage[1891] =  13'b0000000000000; // 0 4.7031538997543976e-05
storage[1892] =  13'b0000100110101; // 309 0.0754273384809494
storage[1893] = -13'b0000001101100; // -108 -0.026484694331884384
storage[1894] =  13'b0000101101000; // 360 0.08799068629741669
storage[1895] =  13'b0001010011110; // 670 0.16362015902996063
storage[1896] = -13'b0000100111000; // -312 -0.07610874623060226
storage[1897] =  13'b0000000000001; // 1 0.00018283944518771023
storage[1898] = -13'b0000011101111; // -239 -0.058405350893735886
storage[1899] = -13'b0000101101101; // -365 -0.08914487063884735
storage[1900] =  13'b0000101011110; // 350 0.08535539358854294
storage[1901] = -13'b0000010111001; // -185 -0.045212700963020325
storage[1902] = -13'b0000011110101; // -245 -0.05985759571194649
storage[1903] = -13'b0000110010011; // -403 -0.09835824370384216
storage[1904] = -13'b0000011100011; // -227 -0.0555235929787159
storage[1905] =  13'b0000011100011; // 227 0.0553734116256237
storage[1906] =  13'b0000010010010; // 146 0.035643767565488815
storage[1907] =  13'b0000010001101; // 141 0.03450499102473259
storage[1908] = -13'b0000001000101; // -69 -0.01678948476910591
storage[1909] = -13'b0000011110001; // -241 -0.05895482748746872
storage[1910] =  13'b0000100110011; // 307 0.07490046322345734
storage[1911] =  13'b0000011010000; // 208 0.05086763948202133
storage[1912] = -13'b0000011101000; // -232 -0.05653905123472214
storage[1913] = -13'b0001001010011; // -595 -0.14520713686943054
storage[1914] = -13'b0000100011101; // -285 -0.06966596096754074
storage[1915] = -13'b0000010011101; // -157 -0.03831082955002785
storage[1916] = -13'b0000101101010; // -362 -0.08846191316843033
storage[1917] = -13'b0000010011000; // -152 -0.03706780821084976
storage[1918] = -13'b0000011111100; // -252 -0.061421871185302734
storage[1919] = -13'b0000010011010; // -154 -0.03766051307320595
storage[1920] = -13'b0000111010001; // -465 -0.11361478269100189
storage[1921] = -13'b0000000101111; // -47 -0.011596065014600754
storage[1922] = -13'b0001000110010; // -562 -0.13731777667999268
storage[1923] = -13'b0000011110000; // -240 -0.058628007769584656
storage[1924] = -13'b0000100010100; // -276 -0.0673411637544632
storage[1925] = -13'b0000100101101; // -301 -0.07345274835824966
storage[1926] =  13'b0000001010001; // 81 0.01986539177596569
storage[1927] =  13'b0001010011100; // 668 0.16319867968559265
storage[1928] =  13'b0000010110100; // 180 0.043868597596883774
storage[1929] = -13'b0000011011010; // -218 -0.05315452441573143
storage[1930] =  13'b0000011100010; // 226 0.05519929528236389
storage[1931] = -13'b0000110001001; // -393 -0.09582588076591492
storage[1932] = -13'b0000001000100; // -68 -0.01654949225485325
storage[1933] = -13'b0000101100000; // -352 -0.0860002264380455
storage[1934] = -13'b0000101100010; // -354 -0.08641863614320755
storage[1935] =  13'b0000101011100; // 348 0.0849483385682106
storage[1936] =  13'b0000000010001; // 17 0.004216640256345272
storage[1937] =  13'b0000000011101; // 29 0.007160961627960205
storage[1938] =  13'b0000100110110; // 310 0.07558383792638779
storage[1939] =  13'b0000110111000; // 440 0.1073286309838295
storage[1940] = -13'b0000000110010; // -50 -0.012203456833958626
storage[1941] =  13'b0000100110111; // 311 0.07596931606531143
storage[1942] =  13'b0001001001010; // 586 0.14299018681049347
storage[1943] =  13'b0000001000101; // 69 0.016837064176797867
storage[1944] =  13'b0000001101111; // 111 0.027010668069124222
storage[1945] =  13'b0000000011010; // 26 0.0064174337312579155
storage[1946] = -13'b0001000011101; // -541 -0.13219007849693298
storage[1947] = -13'b0001000011111; // -543 -0.1325310617685318
storage[1948] =  13'b0000100001000; // 264 0.06452606618404388
storage[1949] = -13'b0000001010011; // -83 -0.020260492339730263
storage[1950] = -13'b0000001001111; // -79 -0.019241992384195328
storage[1951] =  13'b0001010010001; // 657 0.16041885316371918
storage[1952] =  13'b0000110000000; // 384 0.09366375207901001
storage[1953] =  13'b0000010100110; // 166 0.04055342078208923
storage[1954] = -13'b0000000110100; // -52 -0.012684663757681847
storage[1955] =  13'b0000000010011; // 19 0.0046868762001395226
storage[1956] =  13'b0000101100110; // 358 0.08730898797512054
storage[1957] = -13'b0000100110011; // -307 -0.07506230473518372
storage[1958] = -13'b0000110111001; // -441 -0.10766628384590149
storage[1959] =  13'b0000000101100; // 44 0.010745113715529442
storage[1960] =  13'b0000100110100; // 308 0.07510583102703094
storage[1961] = -13'b0000010011011; // -155 -0.03783208876848221
storage[1962] =  13'b0000111111010; // 506 0.12348628789186478
storage[1963] =  13'b0000101010100; // 340 0.0829649269580841
storage[1964] = -13'b0000011111110; // -254 -0.061920758336782455
storage[1965] =  13'b0000101011100; // 348 0.0849713683128357
storage[1966] = -13'b0000000101111; // -47 -0.011423872783780098
storage[1967] = -13'b0000101001100; // -332 -0.08116079121828079
storage[1968] =  13'b0000001100100; // 100 0.024390993639826775
storage[1969] =  13'b0000111100001; // 481 0.1174926683306694
storage[1970] =  13'b0000010100101; // 165 0.04028308019042015
storage[1971] =  13'b0000011110001; // 241 0.05876065418124199
storage[1972] =  13'b0000111010010; // 466 0.11383730173110962
storage[1973] =  13'b0000100110100; // 308 0.07519408315420151
storage[1974] =  13'b0000010110110; // 182 0.04442844167351723
storage[1975] =  13'b0000100110001; // 305 0.0745055228471756
storage[1976] =  13'b0000000100101; // 37 0.008911648765206337
storage[1977] =  13'b0000110100000; // 416 0.10157273709774017
storage[1978] = -13'b0000111011000; // -472 -0.11534490436315536
storage[1979] = -13'b0000111011110; // -478 -0.11674199253320694
storage[1980] =  13'b0000111000101; // 453 0.11070757359266281
storage[1981] =  13'b0000100100111; // 295 0.07204066216945648
storage[1982] = -13'b0000000010011; // -19 -0.004757053218781948
storage[1983] = -13'b0001001000100; // -580 -0.1415734887123108
storage[1984] = -13'b0000001000111; // -71 -0.017455995082855225
storage[1985] = -13'b0000011001011; // -203 -0.049622032791376114
storage[1986] = -13'b0000000101100; // -44 -0.010628740303218365
storage[1987] = -13'b0001001110000; // -624 -0.15237127244472504
storage[1988] = -13'b0001001001010; // -586 -0.14304472506046295
storage[1989] =  13'b0000010101110; // 174 0.04240062087774277
storage[1990] =  13'b0000000101011; // 43 0.010551816783845425
storage[1991] = -13'b0000000111011; // -59 -0.014384971931576729
storage[1992] =  13'b0000000011101; // 29 0.007071352563798428
storage[1993] =  13'b0000100000010; // 258 0.06301604211330414
storage[1994] =  13'b0000010011101; // 157 0.03835981711745262
storage[1995] =  13'b0000101001111; // 335 0.08186770975589752
storage[1996] = -13'b0000011111010; // -250 -0.06108897179365158
storage[1997] = -13'b0000001010101; // -85 -0.02080332115292549
storage[1998] = -13'b0000000000010; // -2 -0.0006001368747092783
storage[1999] = -13'b0000101110100; // -372 -0.09081149846315384
storage[2000] =  13'b0000000011110; // 30 0.007377581670880318
storage[2001] =  13'b0000010101100; // 172 0.041973888874053955
storage[2002] = -13'b0000011011101; // -221 -0.05399394780397415
storage[2003] =  13'b0000100110010; // 306 0.07465535402297974
storage[2004] =  13'b0000001001000; // 72 0.01756509579718113
storage[2005] = -13'b0000100101111; // -303 -0.07399628311395645
storage[2006] = -13'b0000010011001; // -153 -0.03740246593952179
storage[2007] = -13'b0000001001011; // -75 -0.01823147013783455
storage[2008] = -13'b0000010101001; // -169 -0.04114105552434921
storage[2009] = -13'b0000011101100; // -236 -0.05767088755965233
storage[2010] = -13'b0001000111110; // -574 -0.14010176062583923
storage[2011] = -13'b0000100011001; // -281 -0.06867741793394089
storage[2012] =  13'b0000001011011; // 91 0.02217770554125309
storage[2013] =  13'b0000100111010; // 314 0.07672679424285889
storage[2014] = -13'b0000000100110; // -38 -0.009350398555397987
storage[2015] =  13'b0000011111000; // 248 0.06055944412946701
storage[2016] =  13'b0000100011100; // 284 0.06928049772977829
storage[2017] = -13'b0000011011000; // -216 -0.05268684774637222
storage[2018] = -13'b0000000001111; // -15 -0.0036754761822521687
storage[2019] = -13'b0000001110000; // -112 -0.027429824694991112
storage[2020] = -13'b0000000110101; // -53 -0.012873155996203423
storage[2021] = -13'b0001000010100; // -532 -0.12990909814834595
storage[2022] =  13'b0000001110011; // 115 0.02813626080751419
storage[2023] = -13'b0000010011101; // -157 -0.03833361715078354
storage[2024] = -13'b0001010110001; // -689 -0.16831181943416595
storage[2025] = -13'b0000110000010; // -386 -0.09416099637746811
storage[2026] = -13'b0000011011101; // -221 -0.0540202297270298
storage[2027] =  13'b0000010010000; // 144 0.03510028123855591
storage[2028] = -13'b0000010011101; // -157 -0.03833813965320587
storage[2029] =  13'b0000110011110; // 414 0.10114981979131699
storage[2030] =  13'b0000011010001; // 209 0.051086049526929855
storage[2031] = -13'b0000010011001; // -153 -0.03738807141780853
storage[2032] = -13'b0000111000010; // -450 -0.10985727608203888
storage[2033] =  13'b0000001110100; // 116 0.028436115011572838
storage[2034] =  13'b0000100010111; // 279 0.06819544732570648
storage[2035] = -13'b0000111001000; // -456 -0.11121520400047302
storage[2036] = -13'b0000001010011; // -83 -0.020150454714894295
storage[2037] =  13'b0000000101011; // 43 0.010611500591039658
storage[2038] =  13'b0000111100010; // 482 0.117612324655056
storage[2039] =  13'b0000101110010; // 370 0.09026617556810379
storage[2040] =  13'b0000000111001; // 57 0.013945331797003746
storage[2041] =  13'b0000110101011; // 427 0.10420294851064682
storage[2042] =  13'b0000110010000; // 400 0.09766168892383575
storage[2043] =  13'b0000010001101; // 141 0.03430375084280968
storage[2044] =  13'b0000100001110; // 270 0.06598113477230072
storage[2045] = -13'b0000011011101; // -221 -0.053976695984601974
storage[2046] = -13'b0001100100001; // -801 -0.19564814865589142
storage[2047] = -13'b0000011001000; // -200 -0.04877317696809769
storage[2048] = -13'b0001010011001; // -665 -0.16241592168807983
storage[2049] = -13'b0000111101001; // -489 -0.11934619396924973
storage[2050] =  13'b0000000011111; // 31 0.007614989299327135
storage[2051] =  13'b0000100101010; // 298 0.07283302396535873
storage[2052] =  13'b0000100111010; // 314 0.07665538787841797
storage[2053] =  13'b0000110010001; // 401 0.09793484956026077
storage[2054] =  13'b0000011100000; // 224 0.05478533357381821
storage[2055] =  13'b0000000110111; // 55 0.013360939919948578
storage[2056] =  13'b0000010101111; // 175 0.04261818900704384
storage[2057] = -13'b0001010010101; // -661 -0.16148149967193604
storage[2058] = -13'b0010100001111; // -1295 -0.31619223952293396
storage[2059] =  13'b0001000011011; // 539 0.13149797916412354
storage[2060] =  13'b0000001100111; // 103 0.025070933625102043
storage[2061] = -13'b0001000011111; // -543 -0.13252004981040955
storage[2062] =  13'b0001010011110; // 670 0.1635832041501999
storage[2063] =  13'b0000110111111; // 447 0.10918829590082169
storage[2064] = -13'b0000111100001; // -481 -0.11754288524389267
storage[2065] = -13'b0000001001011; // -75 -0.018196599557995796
storage[2066] = -13'b0000000010111; // -23 -0.005600528325885534
storage[2067] = -13'b0000001000111; // -71 -0.017264211550354958
storage[2068] = -13'b0001000000111; // -519 -0.12662017345428467
storage[2069] = -13'b0000000000111; // -7 -0.0016724979504942894
storage[2070] =  13'b0000000010100; // 20 0.0048341648653149605
storage[2071] = -13'b0000001110111; // -119 -0.028992831707000732
storage[2072] = -13'b0000001100001; // -97 -0.023665476590394974
storage[2073] =  13'b0000111101100; // 492 0.12006525695323944
storage[2074] = -13'b0000011100101; // -229 -0.05579269304871559
storage[2075] = -13'b0000001111001; // -121 -0.0295672956854105
storage[2076] =  13'b0000100000010; // 258 0.06310022622346878
storage[2077] = -13'b0000110001110; // -398 -0.09716805070638657
storage[2078] = -13'b0000100101001; // -297 -0.07238879054784775
storage[2079] = -13'b0000001101110; // -110 -0.026774996891617775
storage[2080] =  13'b0000011100000; // 224 0.0547749362885952
storage[2081] =  13'b0000000010101; // 21 0.005206965375691652
storage[2082] =  13'b0000110010011; // 403 0.09839532524347305
storage[2083] =  13'b0000111001110; // 462 0.11275272816419601
storage[2084] = -13'b0000110100010; // -418 -0.10195637494325638
storage[2085] = -13'b0000111110111; // -503 -0.12273012101650238
storage[2086] =  13'b0000010011010; // 154 0.03758516162633896
storage[2087] =  13'b0000011010000; // 208 0.05071501433849335
storage[2088] = -13'b0000100010101; // -277 -0.06768874078989029
storage[2089] = -13'b0000010011100; // -156 -0.03802607208490372
storage[2090] = -13'b0000111000100; // -452 -0.11042635887861252
storage[2091] = -13'b0000110011110; // -414 -0.1011328175663948
storage[2092] =  13'b0000011011010; // 218 0.053225889801979065
storage[2093] = -13'b0000000000001; // -1 -0.0001855501177487895
storage[2094] =  13'b0000010110101; // 181 0.04427528753876686
storage[2095] = -13'b0000010000101; // -133 -0.032565485686063766
storage[2096] = -13'b0000000100011; // -35 -0.008657680824398994
storage[2097] =  13'b0000111100111; // 487 0.11898960173130035
storage[2098] =  13'b0000001100101; // 101 0.02455928735435009
storage[2099] =  13'b0000010111001; // 185 0.045144930481910706
storage[2100] =  13'b0001001110010; // 626 0.15292634069919586
storage[2101] =  13'b0000011011010; // 218 0.05330647528171539
storage[2102] = -13'b0000001000110; // -70 -0.01714520901441574
storage[2103] = -13'b0000100011101; // -285 -0.06953968852758408
storage[2104] = -13'b0000001011110; // -94 -0.022877927869558334
storage[2105] = -13'b0000111011001; // -473 -0.11556325852870941
storage[2106] = -13'b0001011001000; // -712 -0.17373377084732056
storage[2107] =  13'b0000000100001; // 33 0.008046295493841171
storage[2108] = -13'b0001000001000; // -520 -0.12704496085643768
storage[2109] = -13'b0001001100100; // -612 -0.1493503600358963
storage[2110] =  13'b0000010000000; // 128 0.03126435726881027
storage[2111] =  13'b0000110000101; // 389 0.09496182948350906
storage[2112] =  13'b0000001011101; // 93 0.02262810990214348
storage[2113] =  13'b0000001111011; // 123 0.030084148049354553
storage[2114] =  13'b0000100100101; // 293 0.07146509736776352
storage[2115] =  13'b0001001000110; // 582 0.1420809030532837
storage[2116] = -13'b0000001001000; // -72 -0.017686696723103523
storage[2117] =  13'b0000000111001; // 57 0.01398316491395235
storage[2118] =  13'b0000111111000; // 504 0.1230718120932579
storage[2119] = -13'b0001000000111; // -519 -0.12669803202152252
storage[2120] =  13'b0000100011011; // 283 0.06914696097373962
storage[2121] =  13'b0000111101011; // 491 0.1199275553226471
storage[2122] =  13'b0000001110110; // 118 0.02877066656947136
storage[2123] =  13'b0000010000011; // 131 0.03206685930490494
storage[2124] =  13'b0000100000101; // 261 0.06367864459753036
storage[2125] =  13'b0000011000100; // 196 0.04777996614575386
storage[2126] =  13'b0000010101010; // 170 0.04158265143632889
storage[2127] = -13'b0000010101000; // -168 -0.04108817130327225
storage[2128] =  13'b0000001111000; // 120 0.029365038499236107
storage[2129] =  13'b0000100000000; // 256 0.062419045716524124
storage[2130] =  13'b0000100000100; // 260 0.06343933939933777
storage[2131] = -13'b0001100011110; // -798 -0.1947413682937622
storage[2132] =  13'b0000010110011; // 179 0.04364456236362457
storage[2133] = -13'b0001000101110; // -558 -0.13622121512889862
storage[2134] =  13'b0000111100100; // 484 0.11807580292224884
storage[2135] =  13'b0000100011001; // 281 0.06863602995872498
storage[2136] =  13'b0000100111010; // 314 0.07671353220939636
storage[2137] = -13'b0000000111001; // -57 -0.013991528190672398
storage[2138] =  13'b0000110011000; // 408 0.09966319054365158
storage[2139] =  13'b0000010100011; // 163 0.03968055546283722
storage[2140] = -13'b0001001110111; // -631 -0.15396180748939514
storage[2141] =  13'b0000011001000; // 200 0.048777058720588684
storage[2142] =  13'b0000001101101; // 109 0.02673325315117836
storage[2143] =  13'b0000110011010; // 410 0.09999671578407288
storage[2144] =  13'b0000111000101; // 453 0.1105256900191307
storage[2145] = -13'b0000010001001; // -137 -0.03337562084197998
storage[2146] = -13'b0000010100010; // -162 -0.039489347487688065
storage[2147] =  13'b0000110010011; // 403 0.0983872041106224
storage[2148] = -13'b0000000100111; // -39 -0.009414195083081722
storage[2149] =  13'b0000000101101; // 45 0.011075932532548904
storage[2150] =  13'b0000010010011; // 147 0.03598397597670555
storage[2151] =  13'b0000001011011; // 91 0.022135168313980103
storage[2152] =  13'b0000111110110; // 502 0.12254717200994492
storage[2153] = -13'b0000001011011; // -91 -0.02229483611881733
storage[2154] = -13'b0000000000011; // -3 -0.0007814208511263132
storage[2155] = -13'b0001100110110; // -822 -0.20058010518550873
storage[2156] = -13'b0000111001000; // -456 -0.11136018484830856
storage[2157] =  13'b0000100000110; // 262 0.06386714428663254
storage[2158] = -13'b0001100011011; // -795 -0.1941167265176773
storage[2159] = -13'b0000101001101; // -333 -0.08140284568071365
storage[2160] =  13'b0000000000011; // 3 0.0006667338311672211
storage[2161] = -13'b0000000000011; // -3 -0.0006443365127779543
storage[2162] = -13'b0000001010110; // -86 -0.02110472321510315
storage[2163] = -13'b0000000011011; // -27 -0.006525751668959856
storage[2164] = -13'b0000011001100; // -204 -0.04970937967300415
storage[2165] =  13'b0000101001011; // 331 0.080820731818676
storage[2166] =  13'b0000000100101; // 37 0.009079381823539734
storage[2167] = -13'b0000011111101; // -253 -0.06186627969145775
storage[2168] =  13'b0000011011110; // 222 0.054163143038749695
storage[2169] = -13'b0000010111101; // -189 -0.04611770436167717
storage[2170] =  13'b0000011111010; // 250 0.060944825410842896
storage[2171] = -13'b0000000001100; // -12 -0.0030361937824636698
storage[2172] = -13'b0000010011010; // -154 -0.037595234811306
storage[2173] = -13'b0000100111010; // -314 -0.07661660015583038
storage[2174] = -13'b0000101010101; // -341 -0.08319693058729172
storage[2175] = -13'b0000110010100; // -404 -0.0986987054347992
storage[2176] = -13'b0001100000101; // -773 -0.1886059194803238
storage[2177] =  13'b0000100001010; // 266 0.06494330614805222
storage[2178] =  13'b0000011100100; // 228 0.05555685609579086
storage[2179] = -13'b0000100011000; // -280 -0.06845197826623917
storage[2180] = -13'b0000001000100; // -68 -0.016545070335268974
storage[2181] =  13'b0000000100000; // 32 0.007826566696166992
storage[2182] = -13'b0001110101000; // -936 -0.2284042090177536
storage[2183] =  13'b0000001000000; // 64 0.015671273693442345
storage[2184] =  13'b0000010100001; // 161 0.039418645203113556
storage[2185] = -13'b0001110001011; // -907 -0.22137673199176788
storage[2186] =  13'b0000011101110; // 238 0.058076754212379456
storage[2187] =  13'b0000000111010; // 58 0.014101889915764332
storage[2188] = -13'b0000100010010; // -274 -0.06678492575883865
storage[2189] =  13'b0000100101011; // 299 0.0729018822312355
storage[2190] =  13'b0000100100001; // 289 0.07045550644397736
storage[2191] =  13'b0000001110000; // 112 0.027313021942973137
storage[2192] =  13'b0000111001111; // 463 0.11312252283096313
storage[2193] =  13'b0000100000010; // 258 0.06305725127458572
storage[2194] =  13'b0000010010100; // 148 0.036057621240615845
storage[2195] = -13'b0000000011000; // -24 -0.005853986833244562
storage[2196] = -13'b0000100110111; // -311 -0.07588168978691101
storage[2197] =  13'b0000011011011; // 219 0.053448230028152466
storage[2198] =  13'b0000101000000; // 320 0.07817532867193222
storage[2199] = -13'b0000000101101; // -45 -0.011078997515141964
storage[2200] =  13'b0000011000101; // 197 0.04813367500901222
storage[2201] =  13'b0000110110100; // 436 0.10644325613975525
storage[2202] =  13'b0000011100001; // 225 0.054955754429101944
storage[2203] =  13'b0000101100000; // 352 0.08600834012031555
storage[2204] =  13'b0000000101111; // 47 0.01150263287127018
storage[2205] =  13'b0000001100001; // 97 0.023676155135035515
storage[2206] =  13'b0000111010110; // 470 0.11467885226011276
storage[2207] =  13'b0001000010010; // 530 0.1294003576040268
storage[2208] =  13'b0001011101100; // 748 0.1825852245092392
storage[2209] =  13'b0000001000111; // 71 0.017454512417316437
storage[2210] = -13'b0000010011111; // -159 -0.03892119228839874
storage[2211] =  13'b0000001010101; // 85 0.02084525115787983
storage[2212] =  13'b0000011001001; // 201 0.049134448170661926
storage[2213] = -13'b0000110010100; // -404 -0.09871799498796463
storage[2214] =  13'b0000001001111; // 79 0.01931382529437542
storage[2215] =  13'b0000101111010; // 378 0.09227257966995239
storage[2216] =  13'b0000111100111; // 487 0.11898086965084076
storage[2217] =  13'b0000101010010; // 338 0.08254610002040863
storage[2218] = -13'b0001001101001; // -617 -0.15055051445960999
storage[2219] = -13'b0000100001000; // -264 -0.06436076760292053
storage[2220] = -13'b0000111101101; // -493 -0.12047620117664337
storage[2221] =  13'b0000000110000; // 48 0.011640835553407669
storage[2222] = -13'b0000010000111; // -135 -0.03304896503686905
storage[2223] =  13'b0000001011101; // 93 0.022677013650536537
storage[2224] = -13'b0000110010111; // -407 -0.09945415705442429
storage[2225] = -13'b0000110101101; // -429 -0.1047452911734581
storage[2226] = -13'b0000010001010; // -138 -0.03361476585268974
storage[2227] = -13'b0000000110010; // -50 -0.012124523520469666
storage[2228] = -13'b0000001101100; // -108 -0.026349784806370735
storage[2229] =  13'b0000101101010; // 362 0.08837544918060303
storage[2230] =  13'b0000100010011; // 275 0.06704191863536835
storage[2231] = -13'b0000000001001; // -9 -0.00208156555891037
storage[2232] =  13'b0000010011100; // 156 0.03814772516489029
storage[2233] =  13'b0000010111100; // 188 0.045947134494781494
storage[2234] = -13'b0000100011100; // -284 -0.06932726502418518
storage[2235] = -13'b0000000011011; // -27 -0.0065795062109827995
storage[2236] =  13'b0000100011100; // 284 0.069454625248909
storage[2237] =  13'b0000011010001; // 209 0.05110272020101547
storage[2238] =  13'b0000001011001; // 89 0.021700434386730194
storage[2239] = -13'b0000000001011; // -11 -0.002741482574492693
storage[2240] = -13'b0000011110100; // -244 -0.05946660041809082
storage[2241] = -13'b0000011011101; // -221 -0.053842514753341675
storage[2242] = -13'b0000111101110; // -494 -0.12058966606855392
storage[2243] = -13'b0000100010000; // -272 -0.06649424135684967
storage[2244] = -13'b0001100110011; // -819 -0.19984170794487
storage[2245] = -13'b0000011100010; // -226 -0.05512626841664314
storage[2246] =  13'b0000000101110; // 46 0.01119242049753666
storage[2247] = -13'b0000000100011; // -35 -0.00842367671430111
storage[2248] =  13'b0000010110101; // 181 0.04424938187003136
storage[2249] =  13'b0000101110001; // 369 0.09020674973726273
storage[2250] =  13'b0001000001001; // 521 0.12717141211032867
storage[2251] = -13'b0000100111101; // -317 -0.0773790255188942
storage[2252] = -13'b0000011001111; // -207 -0.05052398890256882
storage[2253] = -13'b0000000111100; // -60 -0.014585742726922035
storage[2254] = -13'b0000010011001; // -153 -0.03739055246114731
storage[2255] = -13'b0000110110100; // -436 -0.10639297217130661
storage[2256] = -13'b0000101100001; // -353 -0.08623955398797989
storage[2257] =  13'b0000010110001; // 177 0.04313819482922554
storage[2258] = -13'b0000001100100; // -100 -0.02451406978070736
storage[2259] =  13'b0000010101111; // 175 0.04260547459125519
storage[2260] = -13'b0000001000111; // -71 -0.017266467213630676
storage[2261] = -13'b0000010101110; // -174 -0.04238155484199524
storage[2262] = -13'b0000000001000; // -8 -0.0018998737214133143
storage[2263] = -13'b0000100111110; // -318 -0.07765647768974304
storage[2264] =  13'b0001000010000; // 528 0.128790482878685
storage[2265] =  13'b0000000101110; // 46 0.011164403520524502
storage[2266] =  13'b0000100110011; // 307 0.0749945193529129
storage[2267] =  13'b0001011010011; // 723 0.1765618771314621
storage[2268] =  13'b0000110000010; // 386 0.09417423605918884
storage[2269] = -13'b0000111101101; // -493 -0.12032514065504074
storage[2270] = -13'b0000111110100; // -500 -0.12217836827039719
storage[2271] =  13'b0000000110100; // 52 0.012697387486696243
storage[2272] = -13'b0000110100111; // -423 -0.10330978035926819
storage[2273] =  13'b0000010010011; // 147 0.03599388524889946
storage[2274] =  13'b0000100000111; // 263 0.0641130730509758
storage[2275] =  13'b0000100010101; // 277 0.06773499399423599
storage[2276] =  13'b0000111001011; // 459 0.1120595633983612
storage[2277] = -13'b0000010101001; // -169 -0.041293878108263016
storage[2278] = -13'b0000001010111; // -87 -0.02125890739262104
storage[2279] = -13'b0000101101101; // -365 -0.08907424658536911
storage[2280] = -13'b0000100000111; // -263 -0.06410679221153259
storage[2281] =  13'b0000010010101; // 149 0.03640485554933548
storage[2282] =  13'b0000100110001; // 305 0.07436032593250275
storage[2283] =  13'b0000100101111; // 303 0.07387170195579529
storage[2284] =  13'b0000110000000; // 384 0.0936359316110611
storage[2285] =  13'b0001100011011; // 795 0.19413237273693085
storage[2286] =  13'b0000001100111; // 103 0.025254573673009872
storage[2287] = -13'b0000001101000; // -104 -0.025340668857097626
storage[2288] = -13'b0000111011110; // -478 -0.1166115328669548
storage[2289] = -13'b0011001100011; // -1635 -0.39928609132766724
storage[2290] = -13'b0000101000100; // -324 -0.07898904383182526
storage[2291] = -13'b0001101011000; // -856 -0.2090694159269333
storage[2292] = -13'b0000011110111; // -247 -0.06033569201827049
storage[2293] = -13'b0000110011110; // -414 -0.10112735629081726
storage[2294] = -13'b0000001100000; // -96 -0.023526297882199287
storage[2295] =  13'b0000111011111; // 479 0.11682714521884918
storage[2296] =  13'b0000010001101; // 141 0.03433743491768837
storage[2297] =  13'b0000001111001; // 121 0.029623279348015785
storage[2298] =  13'b0000100000110; // 262 0.06408064067363739
storage[2299] = -13'b0000000011000; // -24 -0.005879594944417477
storage[2300] = -13'b0000000110001; // -49 -0.012017345055937767
storage[2301] =  13'b0000000000110; // 6 0.0015784940915182233
storage[2302] =  13'b0000000101000; // 40 0.009848704561591148
storage[2303] = -13'b0000011011110; // -222 -0.05423952639102936
storage[2304] = -13'b0000011111111; // -255 -0.062284525483846664
storage[2305] =  13'b0000100011000; // 280 0.06833641231060028
storage[2306] =  13'b0000000011010; // 26 0.006250350270420313
storage[2307] =  13'b0000000010110; // 22 0.005453619174659252
storage[2308] =  13'b0000000111001; // 57 0.013902484439313412
storage[2309] =  13'b0000110101011; // 427 0.10429815202951431
storage[2310] = -13'b0000000010100; // -20 -0.004907483700662851
storage[2311] =  13'b0000001101111; // 111 0.02710290066897869
storage[2312] =  13'b0000100101000; // 296 0.07226145267486572
storage[2313] =  13'b0000100001101; // 269 0.06555645167827606
storage[2314] =  13'b0000000010010; // 18 0.004326078575104475
storage[2315] = -13'b0001001000010; // -578 -0.14118991792201996
storage[2316] = -13'b0000010001001; // -137 -0.033441923558712006
storage[2317] = -13'b0000111100000; // -480 -0.11725416779518127
storage[2318] = -13'b0000100011001; // -281 -0.06858669221401215
storage[2319] = -13'b0000010001110; // -142 -0.03455343097448349
storage[2320] = -13'b0000011110011; // -243 -0.059275586158037186
storage[2321] =  13'b0000001011110; // 94 0.022902704775333405
storage[2322] =  13'b0000011010110; // 214 0.05236685276031494
storage[2323] =  13'b0000011000010; // 194 0.04734814167022705
storage[2324] = -13'b0000001110100; // -116 -0.028240090236067772
storage[2325] = -13'b0000101111100; // -380 -0.09289064258337021
storage[2326] = -13'b0000111001000; // -456 -0.1113358587026596
storage[2327] = -13'b0001000001010; // -522 -0.1275414079427719
storage[2328] =  13'b0000000100011; // 35 0.008648463524878025
storage[2329] = -13'b0000001101001; // -105 -0.02575083263218403
storage[2330] = -13'b0000001111101; // -125 -0.030512208119034767
storage[2331] =  13'b0000011111110; // 254 0.062005914747714996
storage[2332] = -13'b0000010100010; // -162 -0.03957662358880043
storage[2333] = -13'b0000110001000; // -392 -0.09572723507881165
storage[2334] =  13'b0000001000000; // 64 0.015571383759379387
storage[2335] =  13'b0000011010101; // 213 0.05197885259985924
storage[2336] =  13'b0000010100011; // 163 0.03979478403925896
storage[2337] =  13'b0000010100110; // 166 0.0405360609292984
storage[2338] =  13'b0000011110000; // 240 0.05858771502971649
storage[2339] =  13'b0000000110010; // 50 0.012319650501012802
storage[2340] = -13'b0000011001100; // -204 -0.04987331107258797
storage[2341] = -13'b0000001010100; // -84 -0.020571043714880943
storage[2342] = -13'b0000110001001; // -393 -0.09583798050880432
storage[2343] = -13'b0001000011001; // -537 -0.13102096319198608
storage[2344] =  13'b0000101101011; // 363 0.08859239518642426
storage[2345] = -13'b0000100101010; // -298 -0.07277841120958328
storage[2346] =  13'b0000000000001; // 1 0.0001890251733129844
storage[2347] = -13'b0000001011010; // -90 -0.021885713562369347
storage[2348] = -13'b0000100010011; // -275 -0.06706058979034424
storage[2349] = -13'b0000011111001; // -249 -0.0608125776052475
storage[2350] = -13'b0001001101000; // -616 -0.15045110881328583
storage[2351] = -13'b0000101110010; // -370 -0.09021258354187012
storage[2352] =  13'b0000001001000; // 72 0.017463715746998787
storage[2353] = -13'b0000011010011; // -211 -0.051436711102724075
storage[2354] = -13'b0000101110011; // -371 -0.09056829661130905
storage[2355] = -13'b0000100011010; // -282 -0.06896859407424927
storage[2356] =  13'b0000001001000; // 72 0.017482463270425797
storage[2357] =  13'b0000110101001; // 425 0.10384505242109299
storage[2358] = -13'b0000000110000; // -48 -0.011800351552665234
storage[2359] = -13'b0000101001001; // -329 -0.08023764938116074
storage[2360] = -13'b0000011100100; // -228 -0.05568030849099159
storage[2361] = -13'b0000010100100; // -164 -0.03999948874115944
storage[2362] = -13'b0000001110001; // -113 -0.027599472552537918
storage[2363] = -13'b0000011110110; // -246 -0.06009995937347412
storage[2364] = -13'b0000001111011; // -123 -0.029979011043906212
storage[2365] = -13'b0000011001011; // -203 -0.04944460466504097
storage[2366] = -13'b0000110110000; // -432 -0.10535703599452972
storage[2367] = -13'b0000100000110; // -262 -0.06385128200054169
storage[2368] =  13'b0000001100011; // 99 0.024231506511569023
storage[2369] =  13'b0000011101101; // 237 0.05783016234636307
storage[2370] =  13'b0000101010000; // 336 0.08203639090061188
storage[2371] = -13'b0000001001000; // -72 -0.01754802279174328
storage[2372] =  13'b0000001011011; // 91 0.022122304886579514
storage[2373] =  13'b0001010010011; // 659 0.16080909967422485
storage[2374] = -13'b0000010010000; // -144 -0.0350443497300148
storage[2375] = -13'b0000011110000; // -240 -0.058603305369615555
storage[2376] = -13'b0000011001001; // -201 -0.04915396124124527
storage[2377] =  13'b0001010110000; // 688 0.16804876923561096
storage[2378] =  13'b0000101101001; // 361 0.08822233229875565
storage[2379] =  13'b0000101110010; // 370 0.09043542295694351
storage[2380] =  13'b0000100010010; // 274 0.06701555103063583
storage[2381] = -13'b0000010110011; // -179 -0.04369862377643585
storage[2382] = -13'b0000000100010; // -34 -0.008290656842291355
storage[2383] =  13'b0000000001101; // 13 0.003264929633587599
storage[2384] =  13'b0000001010110; // 86 0.02099551260471344
storage[2385] = -13'b0000010000100; // -132 -0.03214545175433159
storage[2386] = -13'b0000111001100; // -460 -0.11237943172454834
storage[2387] = -13'b0000010101010; // -170 -0.041520729660987854
storage[2388] = -13'b0000000010010; // -18 -0.004366767592728138
storage[2389] = -13'b0000010011100; // -156 -0.03814135864377022
storage[2390] = -13'b0000000000011; // -3 -0.0007485761307179928
storage[2391] = -13'b0000000100101; // -37 -0.009096070192754269
storage[2392] =  13'b0000001011111; // 95 0.023157551884651184
storage[2393] =  13'b0000010010010; // 146 0.03557996824383736
storage[2394] =  13'b0000010111111; // 191 0.04653483256697655
storage[2395] = -13'b0001001111110; // -638 -0.15564242005348206
storage[2396] = -13'b0000010110000; // -176 -0.04307137429714203
storage[2397] =  13'b0000011110001; // 241 0.058912813663482666
storage[2398] = -13'b0000010010010; // -146 -0.035559702664613724
storage[2399] =  13'b0000100010001; // 273 0.06671546399593353
storage[2400] =  13'b0000010110110; // 182 0.04446117952466011
storage[2401] =  13'b0000100011110; // 286 0.06974294781684875
storage[2402] =  13'b0000110101101; // 429 0.10484527051448822
storage[2403] =  13'b0000010011011; // 155 0.03779733180999756
storage[2404] = -13'b0000111001101; // -461 -0.1126386821269989
storage[2405] = -13'b0000011001000; // -200 -0.04892803728580475
storage[2406] =  13'b0000000111101; // 61 0.014773777686059475
storage[2407] = -13'b0000101111101; // -381 -0.09311174601316452
storage[2408] =  13'b0000001001011; // 75 0.018371980637311935
storage[2409] = -13'b0000001001000; // -72 -0.017557531595230103
storage[2410] = -13'b0000111000011; // -451 -0.11015024781227112
storage[2411] =  13'b0000010000110; // 134 0.03274095803499222
storage[2412] =  13'b0000000010100; // 20 0.004857651423662901
storage[2413] = -13'b0001010110101; // -693 -0.16930752992630005
storage[2414] = -13'b0010110111111; // -1471 -0.3591171205043793
storage[2415] = -13'b0001010011111; // -671 -0.16374512016773224
storage[2416] = -13'b0010010100101; // -1189 -0.29022809863090515
storage[2417] = -13'b0001101111001; // -889 -0.21692368388175964
storage[2418] = -13'b0000011100001; // -225 -0.054931122809648514
storage[2419] = -13'b0001101101010; // -874 -0.21328456699848175
storage[2420] = -13'b0000010111100; // -188 -0.04600181430578232
storage[2421] =  13'b0000001001101; // 77 0.01879044435918331
storage[2422] =  13'b0000100111010; // 314 0.07668720185756683
storage[2423] = -13'b0000100011000; // -280 -0.06839026510715485
storage[2424] =  13'b0000101111011; // 379 0.09255574643611908
storage[2425] =  13'b0000001011000; // 88 0.02151375636458397
storage[2426] = -13'b0000000101001; // -41 -0.009934010915458202
storage[2427] =  13'b0000000001100; // 12 0.002957841381430626
storage[2428] = -13'b0000001101111; // -111 -0.027098486199975014
storage[2429] = -13'b0000000111111; // -63 -0.015386605635285378
storage[2430] =  13'b0000010111100; // 188 0.04596952348947525
storage[2431] =  13'b0000100110100; // 308 0.07514090836048126
storage[2432] =  13'b0000100100100; // 292 0.0713726207613945
storage[2433] =  13'b0000001010110; // 86 0.020974496379494667
storage[2434] =  13'b0000011101101; // 237 0.05794860050082207
storage[2435] =  13'b0000010101111; // 175 0.04268302768468857
storage[2436] = -13'b0000001011101; // -93 -0.022623741999268532
storage[2437] = -13'b0000001111111; // -127 -0.030943894758820534
storage[2438] =  13'b0000111101001; // 489 0.11945280432701111
storage[2439] =  13'b0000011000010; // 194 0.04747087135910988
storage[2440] = -13'b0000100110100; // -308 -0.07530876249074936
storage[2441] = -13'b0001101101000; // -872 -0.21299780905246735
storage[2442] = -13'b0010001111111; // -1151 -0.28102555871009827
storage[2443] = -13'b0000110000011; // -387 -0.09460004419088364
storage[2444] = -13'b0000001110111; // -119 -0.029060116037726402
storage[2445] =  13'b0000000110101; // 53 0.0128253772854805
storage[2446] =  13'b0000100010001; // 273 0.06661329418420792
storage[2447] =  13'b0000100011101; // 285 0.06955164670944214
storage[2448] =  13'b0000000110101; // 53 0.013016795739531517
storage[2449] =  13'b0000000100110; // 38 0.009282216429710388
storage[2450] =  13'b0000001000000; // 64 0.015508373267948627
storage[2451] =  13'b0000110111001; // 441 0.10773272067308426
storage[2452] =  13'b0000110010111; // 407 0.09935963898897171
storage[2453] =  13'b0000011101010; // 234 0.05713873729109764
storage[2454] =  13'b0000001010000; // 80 0.01961429975926876
storage[2455] =  13'b0000101000001; // 321 0.07826214283704758
storage[2456] =  13'b0001001010011; // 595 0.14527590572834015
storage[2457] =  13'b0000010001111; // 143 0.034963835030794144
storage[2458] = -13'b0000100001110; // -270 -0.06593920290470123
storage[2459] = -13'b0000101010011; // -339 -0.08269311487674713
storage[2460] = -13'b0000101100101; // -357 -0.08713436126708984
storage[2461] = -13'b0000110001010; // -394 -0.096165232360363
storage[2462] =  13'b0000001100011; // 99 0.024106059223413467
storage[2463] = -13'b0000001100000; // -96 -0.02350415661931038
storage[2464] =  13'b0000011001000; // 200 0.048729002475738525
storage[2465] =  13'b0000001001011; // 75 0.01841200888156891
storage[2466] =  13'b0000100100100; // 292 0.07129693031311035
storage[2467] =  13'b0000100110000; // 304 0.07411517202854156
storage[2468] =  13'b0000000010000; // 16 0.003786020912230015
storage[2469] =  13'b0000010111010; // 186 0.04551176726818085
storage[2470] = -13'b0000010011000; // -152 -0.03719491511583328
storage[2471] = -13'b0000010100011; // -163 -0.03969281166791916
storage[2472] = -13'b0000011010111; // -215 -0.052435439079999924
storage[2473] =  13'b0000010010010; // 146 0.03555485978722572
storage[2474] =  13'b0000101101101; // 365 0.08904582262039185
storage[2475] =  13'b0000100111111; // 319 0.07787437736988068
storage[2476] = -13'b0000000000111; // -7 -0.001607144600711763
storage[2477] = -13'b0000000000001; // -1 -0.0003194813907612115
storage[2478] =  13'b0000001001100; // 76 0.018589885905385017
storage[2479] =  13'b0000011001111; // 207 0.05065853148698807
storage[2480] =  13'b0000000110000; // 48 0.011694776825606823
storage[2481] = -13'b0000111001000; // -456 -0.11137772351503372
storage[2482] =  13'b0000001101100; // 108 0.02629907801747322
storage[2483] = -13'b0000110010101; // -405 -0.09880269318819046
storage[2484] = -13'b0001111010000; // -976 -0.23831775784492493
storage[2485] = -13'b0000010000101; // -133 -0.0324445441365242
storage[2486] = -13'b0000000110101; // -53 -0.013044847175478935
storage[2487] =  13'b0000101000011; // 323 0.07886449247598648
storage[2488] = -13'b0000101110101; // -373 -0.09113849699497223
storage[2489] =  13'b0000001110100; // 116 0.028396278619766235
storage[2490] =  13'b0000111110001; // 497 0.12144049257040024
storage[2491] =  13'b0001010110101; // 693 0.16911546885967255
storage[2492] = -13'b0000111001101; // -461 -0.11261912435293198
storage[2493] = -13'b0000100011000; // -280 -0.06824960559606552
storage[2494] =  13'b0000001011011; // 91 0.02219310961663723
storage[2495] =  13'b0000010011101; // 157 0.038431014865636826
storage[2496] = -13'b0000000010010; // -18 -0.004331725183874369
storage[2497] = -13'b0000010000011; // -131 -0.032083719968795776
storage[2498] = -13'b0000001001101; // -77 -0.018731527030467987
storage[2499] = -13'b0000011101011; // -235 -0.05728224292397499
storage[2500] =  13'b0001010010111; // 663 0.16190288960933685
storage[2501] =  13'b0000110011001; // 409 0.09992853552103043
storage[2502] = -13'b0000100001010; // -266 -0.06489484757184982
storage[2503] =  13'b0000100010101; // 277 0.06758267432451248
storage[2504] =  13'b0000010100000; // 160 0.03896259143948555
storage[2505] = -13'b0000001100011; // -99 -0.024174172431230545
storage[2506] = -13'b0000000010100; // -20 -0.0048821973614394665
storage[2507] = -13'b0000100111110; // -318 -0.07754026353359222
storage[2508] = -13'b0000000110011; // -51 -0.012333212420344353
storage[2509] =  13'b0000010010100; // 148 0.0362243726849556
storage[2510] = -13'b0000000011101; // -29 -0.007002802565693855
storage[2511] = -13'b0000001100001; // -97 -0.02357739396393299
storage[2512] =  13'b0000010000001; // 129 0.0315316841006279
storage[2513] =  13'b0000001101001; // 105 0.025680629536509514
storage[2514] =  13'b0000010011100; // 156 0.03816094622015953
storage[2515] = -13'b0000010011100; // -156 -0.03807641938328743
storage[2516] =  13'b0000000001000; // 8 0.0019740310963243246
storage[2517] =  13'b0000010000010; // 130 0.03175684064626694
storage[2518] = -13'b0000110000101; // -389 -0.09492567181587219
storage[2519] = -13'b0000100100111; // -295 -0.07208354026079178
storage[2520] =  13'b0000001001011; // 75 0.018420755863189697
storage[2521] = -13'b0000000001100; // -12 -0.0029391988646239042
storage[2522] = -13'b0000000001100; // -12 -0.003048934042453766
storage[2523] = -13'b0000001101111; // -111 -0.02718968503177166
storage[2524] = -13'b0000011011010; // -218 -0.05330273509025574
storage[2525] = -13'b0001001111111; // -639 -0.15603835880756378
storage[2526] = -13'b0001100100001; // -801 -0.19564634561538696
storage[2527] =  13'b0000100010011; // 275 0.06719741225242615
storage[2528] = -13'b0000000111000; // -56 -0.013599221594631672
storage[2529] = -13'b0000011010110; // -214 -0.05229712650179863
storage[2530] = -13'b0000000110000; // -48 -0.01173901092261076
storage[2531] = -13'b0000010110100; // -180 -0.043957244604825974
storage[2532] = -13'b0000001101011; // -107 -0.026005765423178673
storage[2533] = -13'b0000010010010; // -146 -0.03561649098992348
storage[2534] =  13'b0000111011101; // 477 0.11655936390161514
storage[2535] =  13'b0001100001000; // 776 0.18934659659862518
storage[2536] =  13'b0000111111001; // 505 0.12326869368553162
storage[2537] =  13'b0000101110011; // 371 0.09061674028635025
storage[2538] =  13'b0000011110100; // 244 0.059526778757572174
storage[2539] =  13'b0000001101101; // 109 0.026670895516872406
storage[2540] =  13'b0000010011000; // 152 0.03710814192891121
storage[2541] = -13'b0000000011100; // -28 -0.006948643364012241
storage[2542] =  13'b0000010011010; // 154 0.037643738090991974
storage[2543] =  13'b0000100100000; // 288 0.07036518305540085
storage[2544] =  13'b0000000000000; // 0 2.302958455402404e-05
storage[2545] =  13'b0000000001110; // 14 0.003461417043581605
storage[2546] =  13'b0000011110011; // 243 0.0594334676861763
storage[2547] =  13'b0000010111011; // 187 0.04575758054852486
storage[2548] = -13'b0000000100001; // -33 -0.00810952391475439
storage[2549] =  13'b0000001110001; // 113 0.02752692997455597
storage[2550] =  13'b0000100101011; // 299 0.07296708971261978
storage[2551] = -13'b0000010001101; // -141 -0.03444085642695427
storage[2552] = -13'b0000011110111; // -247 -0.06035977974534035
storage[2553] =  13'b0000011111111; // 255 0.06233514845371246
storage[2554] = -13'b0000000110000; // -48 -0.011692616157233715
storage[2555] =  13'b0000000000011; // 3 0.0007078346097841859
storage[2556] =  13'b0001000001110; // 526 0.12842223048210144
storage[2557] =  13'b0000100100010; // 290 0.07074832171201706
storage[2558] =  13'b0001000011011; // 539 0.13150466978549957
storage[2559] =  13'b0000001010010; // 82 0.020014720037579536
storage[2560] =  13'b0000000010011; // 19 0.004662424325942993
storage[2561] =  13'b0001000010101; // 533 0.13002772629261017
storage[2562] = -13'b0000011011010; // -218 -0.0532265305519104
storage[2563] =  13'b0000010111100; // 188 0.04579586535692215
storage[2564] =  13'b0001011110000; // 752 0.18362411856651306
storage[2565] =  13'b0000010111011; // 187 0.04571985453367233
storage[2566] =  13'b0001001111011; // 635 0.15507858991622925
storage[2567] = -13'b0001010011011; // -667 -0.1628996878862381
storage[2568] = -13'b0000100100101; // -293 -0.07160770148038864
storage[2569] = -13'b0000000010110; // -22 -0.00546081131324172
storage[2570] = -13'b0000110010010; // -402 -0.09824805706739426
storage[2571] = -13'b0000001000110; // -70 -0.017194341868162155
storage[2572] =  13'b0000010010100; // 148 0.036089569330215454
storage[2573] =  13'b0000011000100; // 196 0.047860387712717056
storage[2574] =  13'b0000001001011; // 75 0.01835072971880436
storage[2575] =  13'b0000000010011; // 19 0.004748606588691473
storage[2576] =  13'b0000001110000; // 112 0.02723902091383934
storage[2577] = -13'b0000001011110; // -94 -0.022880518808960915
storage[2578] =  13'b0000001111000; // 120 0.029182953760027885
storage[2579] = -13'b0000000011101; // -29 -0.0069630383513867855
storage[2580] = -13'b0000101100010; // -354 -0.08631295710802078
storage[2581] =  13'b0000011000011; // 195 0.047702230513095856
storage[2582] = -13'b0000000101011; // -43 -0.010548458434641361
storage[2583] = -13'b0000001000001; // -65 -0.01597975566983223
storage[2584] =  13'b0000001111001; // 121 0.02954910136759281
storage[2585] =  13'b0000100010100; // 276 0.06728491187095642
storage[2586] =  13'b0000010011011; // 155 0.037747640162706375
storage[2587] =  13'b0000000110100; // 52 0.012760455720126629
storage[2588] =  13'b0000000011101; // 29 0.007036565337330103
storage[2589] =  13'b0000000101100; // 44 0.010679639875888824
storage[2590] = -13'b0000011001100; // -204 -0.04970784857869148
storage[2591] =  13'b0000011000100; // 196 0.04795714095234871
storage[2592] =  13'b0000011010000; // 208 0.0508563369512558
storage[2593] = -13'b0000011110110; // -246 -0.060113321989774704
storage[2594] = -13'b0000110000110; // -390 -0.09517737478017807
storage[2595] = -13'b0000000001000; // -8 -0.001981880748644471
storage[2596] = -13'b0000011101110; // -238 -0.05804469808936119
storage[2597] = -13'b0001010111111; // -703 -0.17154543101787567
storage[2598] = -13'b0000110101000; // -424 -0.10356422513723373
storage[2599] = -13'b0000100100001; // -289 -0.07053888589143753
storage[2600] = -13'b0000011101000; // -232 -0.056740839034318924
storage[2601] =  13'b0000010011110; // 158 0.03846661001443863
storage[2602] =  13'b0000100010011; // 275 0.06725896894931793
storage[2603] =  13'b0000011001110; // 206 0.050369445234537125
storage[2604] = -13'b0000011100000; // -224 -0.0548073872923851
storage[2605] =  13'b0000010011010; // 154 0.037579674273729324
storage[2606] =  13'b0000100000100; // 260 0.06351068615913391
storage[2607] = -13'b0000011000011; // -195 -0.047604598104953766
storage[2608] = -13'b0000000101101; // -45 -0.011069739237427711
storage[2609] =  13'b0000000011000; // 24 0.005864646285772324
storage[2610] =  13'b0000000011000; // 24 0.005865638609975576
storage[2611] =  13'b0000000100111; // 39 0.009489907883107662
storage[2612] =  13'b0000000011010; // 26 0.006356647703796625
storage[2613] =  13'b0001000100101; // 549 0.1339770406484604
storage[2614] = -13'b0000100010111; // -279 -0.0679967850446701
storage[2615] = -13'b0000001110101; // -117 -0.02848251350224018
storage[2616] =  13'b0000100011100; // 284 0.06931211799383163
storage[2617] =  13'b0001000100011; // 547 0.13343806564807892
storage[2618] =  13'b0000010100010; // 162 0.03961217403411865
storage[2619] = -13'b0000001001000; // -72 -0.01750185340642929
storage[2620] = -13'b0000101101101; // -365 -0.08903103321790695
storage[2621] = -13'b0000001111010; // -122 -0.02978093922138214
storage[2622] =  13'b0000011111010; // 250 0.06098199263215065
storage[2623] =  13'b0000101011111; // 351 0.08557768911123276
storage[2624] = -13'b0000110111011; // -443 -0.10819444060325623
storage[2625] = -13'b0001000001111; // -527 -0.12864865362644196
storage[2626] =  13'b0000011001010; // 202 0.04934835806488991
storage[2627] = -13'b0000101000111; // -327 -0.07981516420841217
storage[2628] =  13'b0000011011100; // 220 0.053651317954063416
storage[2629] = -13'b0000111011001; // -473 -0.11552482843399048
storage[2630] = -13'b0000101100110; // -358 -0.08742208778858185
storage[2631] =  13'b0000001001011; // 75 0.018256476148962975
storage[2632] =  13'b0000010001010; // 138 0.03362515568733215
storage[2633] = -13'b0000001100111; // -103 -0.025091305375099182
storage[2634] = -13'b0000101110000; // -368 -0.08991780877113342
storage[2635] =  13'b0000000010000; // 16 0.003926498349756002
storage[2636] = -13'b0000101001010; // -330 -0.08046070486307144
storage[2637] = -13'b0000010110000; // -176 -0.043021898716688156
storage[2638] = -13'b0000010101001; // -169 -0.041267234832048416
storage[2639] = -13'b0000001010000; // -80 -0.01941806636750698
storage[2640] = -13'b0000011101100; // -236 -0.05764824524521828
storage[2641] =  13'b0000111001100; // 460 0.1122300922870636
storage[2642] =  13'b0000011101011; // 235 0.05740957707166672
storage[2643] = -13'b0000010100110; // -166 -0.0404505729675293
storage[2644] =  13'b0001011010010; // 722 0.17619448900222778
storage[2645] =  13'b0001000001011; // 523 0.1276571899652481
storage[2646] = -13'b0000000001000; // -8 -0.0019820339512079954
storage[2647] = -13'b0001001001100; // -588 -0.14354468882083893
storage[2648] = -13'b0000111100100; // -484 -0.11804984509944916
storage[2649] =  13'b0000101010010; // 338 0.08263322710990906
storage[2650] =  13'b0000001010010; // 82 0.019904235377907753
storage[2651] = -13'b0000000101000; // -40 -0.009693105705082417
storage[2652] = -13'b0000000101100; // -44 -0.010687917470932007
storage[2653] =  13'b0001011000100; // 708 0.17295873165130615
storage[2654] =  13'b0000101111000; // 376 0.0919124037027359
storage[2655] = -13'b0000011001000; // -200 -0.04877091571688652
storage[2656] = -13'b0000010100101; // -165 -0.040179431438446045
storage[2657] = -13'b0000000000011; // -3 -0.0006395389791578054
storage[2658] =  13'b0000101001010; // 330 0.08049938082695007
storage[2659] =  13'b0000011001110; // 206 0.05034615099430084
storage[2660] =  13'b0000011011101; // 221 0.05395616590976715
storage[2661] =  13'b0000101000001; // 321 0.07827574014663696
storage[2662] = -13'b0000100011001; // -281 -0.06855497509241104
storage[2663] = -13'b0000001110000; // -112 -0.02726569212973118
storage[2664] = -13'b0000001110000; // -112 -0.02723190002143383
storage[2665] =  13'b0000100110001; // 305 0.07443711906671524
storage[2666] = -13'b0000100101001; // -297 -0.07242385298013687
storage[2667] = -13'b0000101010011; // -339 -0.08279833942651749
storage[2668] =  13'b0001000010000; // 528 0.12891383469104767
storage[2669] = -13'b0000001000100; // -68 -0.01656714454293251
storage[2670] = -13'b0000110110101; // -437 -0.10658891499042511
storage[2671] =  13'b0000101001011; // 331 0.08078128844499588
storage[2672] =  13'b0000010100100; // 164 0.03999588266015053
storage[2673] =  13'b0000110111111; // 447 0.10905895382165909
storage[2674] = -13'b0000010011101; // -157 -0.03834730014204979
storage[2675] = -13'b0000001011111; // -95 -0.02312472090125084
storage[2676] =  13'b0000011111111; // 255 0.062276147305965424
storage[2677] = -13'b0000101010100; // -340 -0.08296220004558563
storage[2678] =  13'b0000010010001; // 145 0.035457316786050797
storage[2679] =  13'b0000011111111; // 255 0.06218218430876732
storage[2680] =  13'b0000100101111; // 303 0.0740724429488182
storage[2681] = -13'b0000100000010; // -258 -0.06297695636749268
storage[2682] = -13'b0000011000001; // -193 -0.04703253135085106
storage[2683] = -13'b0000010001001; // -137 -0.03344608098268509
storage[2684] = -13'b0000001100111; // -103 -0.025188297033309937
storage[2685] =  13'b0000001010001; // 81 0.01970069482922554
storage[2686] =  13'b0000000001000; // 8 0.001912159495986998
storage[2687] = -13'b0000011000111; // -199 -0.048462942242622375
storage[2688] = -13'b0001000100100; // -548 -0.13381415605545044
storage[2689] =  13'b0000100111011; // 315 0.07686813920736313
storage[2690] =  13'b0000100000001; // 257 0.0628332644701004
storage[2691] =  13'b0001001000001; // 577 0.14098024368286133
storage[2692] =  13'b0000000000100; // 4 0.0009301829850301147
storage[2693] = -13'b0000101101000; // -360 -0.08781873434782028
storage[2694] = -13'b0000001111100; // -124 -0.030164914205670357
storage[2695] =  13'b0000111000000; // 448 0.10946142673492432
storage[2696] = -13'b0000010110011; // -179 -0.04373981058597565
storage[2697] =  13'b0000101111111; // 383 0.09355586022138596
storage[2698] = -13'b0001000011100; // -540 -0.13185055553913116
storage[2699] = -13'b0000010111101; // -189 -0.04618668556213379
storage[2700] =  13'b0000000101110; // 46 0.01116659864783287
storage[2701] =  13'b0000000111110; // 62 0.015245688147842884
storage[2702] =  13'b0000010011111; // 159 0.03875422477722168
storage[2703] =  13'b0000000111110; // 62 0.015106319449841976
storage[2704] =  13'b0001001110100; // 628 0.15324321389198303
storage[2705] = -13'b0000001000111; // -71 -0.017286887392401695
storage[2706] =  13'b0000101100001; // 353 0.08623026311397552
storage[2707] = -13'b0000001100111; // -103 -0.025141164660453796
storage[2708] =  13'b0000001010000; // 80 0.019504576921463013
storage[2709] =  13'b0000011101011; // 235 0.057326946407556534
storage[2710] =  13'b0000101110001; // 369 0.09018352627754211
storage[2711] = -13'b0000001100001; // -97 -0.023782650008797646
storage[2712] = -13'b0000011100101; // -229 -0.05592027306556702
storage[2713] =  13'b0000101110111; // 375 0.09152808040380478
storage[2714] = -13'b0000100110000; // -304 -0.07418347150087357
storage[2715] =  13'b0000011011100; // 220 0.05370696261525154
storage[2716] =  13'b0000100011100; // 284 0.06941723823547363
storage[2717] =  13'b0000000011011; // 27 0.0066297403536736965
storage[2718] =  13'b0000111000011; // 451 0.11022664606571198
storage[2719] = -13'b0001000100110; // -550 -0.1343858242034912
storage[2720] = -13'b0000101111110; // -382 -0.09324432909488678
storage[2721] = -13'b0000011000111; // -199 -0.04849938675761223
storage[2722] = -13'b0000110011001; // -409 -0.0998363196849823
storage[2723] = -13'b0001001100111; // -615 -0.15013156831264496
storage[2724] = -13'b0000010101011; // -171 -0.041739460080862045
storage[2725] = -13'b0000100000000; // -256 -0.062418609857559204
storage[2726] = -13'b0000101010010; // -338 -0.08263465017080307
storage[2727] =  13'b0000010100111; // 167 0.04081668704748154
storage[2728] = -13'b0000000010101; // -21 -0.005073670297861099
storage[2729] =  13'b0000110010100; // 404 0.09861022979021072
storage[2730] =  13'b0000000010101; // 21 0.00517334695905447
storage[2731] =  13'b0000000101101; // 45 0.010929100215435028
storage[2732] = -13'b0000100111110; // -318 -0.07770898938179016
storage[2733] = -13'b0000011000010; // -194 -0.04727660492062569
storage[2734] =  13'b0001010010011; // 659 0.16096548736095428
storage[2735] =  13'b0001000111101; // 573 0.1398402601480484
storage[2736] =  13'b0000100110110; // 310 0.07559303194284439
storage[2737] = -13'b0000011110000; // -240 -0.05863180011510849
storage[2738] = -13'b0000010001100; // -140 -0.03420913591980934
storage[2739] = -13'b0000000111001; // -57 -0.01397673599421978
storage[2740] = -13'b0000000011100; // -28 -0.006880135275423527
storage[2741] = -13'b0000011001000; // -200 -0.04878313094377518
storage[2742] =  13'b0000000110000; // 48 0.01179785281419754
storage[2743] = -13'b0000011100001; // -225 -0.05490008741617203
storage[2744] = -13'b0000100011010; // -282 -0.06877806037664413
storage[2745] =  13'b0000000001110; // 14 0.0034414564725011587
storage[2746] = -13'b0000001010110; // -86 -0.020887130871415138
storage[2747] =  13'b0000011110100; // 244 0.05951179563999176
storage[2748] =  13'b0000010101011; // 171 0.04173007234930992
storage[2749] =  13'b0000101100010; // 354 0.08652844280004501
storage[2750] = -13'b0000010000100; // -132 -0.03215542808175087
storage[2751] = -13'b0000100100010; // -290 -0.07072142511606216
storage[2752] =  13'b0000010000100; // 132 0.0322762131690979
storage[2753] =  13'b0000100101011; // 299 0.07304666191339493
storage[2754] =  13'b0000001011001; // 89 0.021705295890569687
storage[2755] = -13'b0000001101011; // -107 -0.026229247450828552
storage[2756] = -13'b0000001100010; // -98 -0.024034319445490837
storage[2757] = -13'b0000001110110; // -118 -0.02876693569123745
storage[2758] =  13'b0000001111010; // 122 0.029734469950199127
storage[2759] =  13'b0000001101110; // 110 0.026772381737828255
storage[2760] = -13'b0000001000111; // -71 -0.01738513447344303
storage[2761] =  13'b0001000101110; // 558 0.13633637130260468
storage[2762] =  13'b0000011001101; // 205 0.05005413293838501
storage[2763] = -13'b0000001111001; // -121 -0.02943389117717743
storage[2764] =  13'b0000000110010; // 50 0.012245703488588333
storage[2765] = -13'b0000010010100; // -148 -0.03621033951640129
storage[2766] = -13'b0000100010101; // -277 -0.067709781229496
storage[2767] =  13'b0000000101101; // 45 0.0109056131914258
storage[2768] =  13'b0001010111100; // 700 0.1708197444677353
storage[2769] =  13'b0000110001011; // 395 0.09647803753614426
storage[2770] =  13'b0000010011000; // 152 0.03716326132416725
storage[2771] =  13'b0001010101001; // 681 0.166183739900589
storage[2772] =  13'b0000000110001; // 49 0.011908076703548431
storage[2773] =  13'b0000001110100; // 116 0.02843024954199791
storage[2774] =  13'b0000000101111; // 47 0.01152388658374548
storage[2775] = -13'b0000000011000; // -24 -0.005778581835329533
storage[2776] =  13'b0000001101000; // 104 0.025345301255583763
storage[2777] =  13'b0000010110010; // 178 0.043550994247198105
storage[2778] = -13'b0000000100101; // -37 -0.008934308774769306
storage[2779] =  13'b0001000100000; // 544 0.1327151358127594
storage[2780] =  13'b0001010010010; // 658 0.1606091856956482
storage[2781] =  13'b0000000001010; // 10 0.00243525137193501
storage[2782] =  13'b0000001010111; // 87 0.021170729771256447
storage[2783] =  13'b0000000111010; // 58 0.014139449223876
storage[2784] = -13'b0000000101010; // -42 -0.010147439315915108
storage[2785] = -13'b0000110111001; // -441 -0.10761963576078415
storage[2786] = -13'b0000000010100; // -20 -0.00486000394448638
storage[2787] =  13'b0000101100011; // 355 0.08655048161745071
storage[2788] =  13'b0000000010111; // 23 0.005534650757908821
storage[2789] =  13'b0000101011001; // 345 0.08427347242832184
storage[2790] =  13'b0000100010101; // 277 0.0676783099770546
storage[2791] = -13'b0000100101011; // -299 -0.07294196635484695
storage[2792] = -13'b0000000110100; // -52 -0.012743971310555935
storage[2793] = -13'b0001000100010; // -546 -0.13340304791927338
storage[2794] = -13'b0000101001000; // -328 -0.07997403293848038
storage[2795] = -13'b0000011011111; // -223 -0.054538339376449585
storage[2796] = -13'b0000001000001; // -65 -0.015834622085094452
storage[2797] =  13'b0000000101010; // 42 0.010260041803121567
storage[2798] =  13'b0000001111110; // 126 0.03070070408284664
storage[2799] =  13'b0000000000100; // 4 0.0010389800881966949
storage[2800] = -13'b0000000110111; // -55 -0.013347042724490166
storage[2801] =  13'b0000010001001; // 137 0.033400628715753555
storage[2802] =  13'b0000001100011; // 99 0.024213038384914398
storage[2803] =  13'b0000101100000; // 352 0.08600980043411255
storage[2804] = -13'b0000000101001; // -41 -0.009978920221328735
storage[2805] = -13'b0000001101111; // -111 -0.027138743549585342
storage[2806] =  13'b0000011111101; // 253 0.061846256256103516
storage[2807] = -13'b0000001001110; // -78 -0.01913209818303585
storage[2808] = -13'b0001000001111; // -527 -0.12873561680316925
storage[2809] = -13'b0000000101000; // -40 -0.00976224523037672
storage[2810] = -13'b0000000100001; // -33 -0.008074592798948288
storage[2811] =  13'b0000000011000; // 24 0.005856725387275219
storage[2812] = -13'b0000100110011; // -307 -0.07489927113056183
storage[2813] = -13'b0000100011010; // -282 -0.06888795644044876
storage[2814] = -13'b0000010110100; // -180 -0.044041454792022705
storage[2815] =  13'b0000001110010; // 114 0.02774965949356556
storage[2816] =  13'b0000010000000; // 128 0.031191295012831688
storage[2817] = -13'b0000001000011; // -67 -0.016321973875164986
storage[2818] =  13'b0000011101110; // 238 0.05800396576523781
storage[2819] = -13'b0000001000001; // -65 -0.015969088301062584
storage[2820] = -13'b0000001110111; // -119 -0.02893466129899025
storage[2821] = -13'b0000011110010; // -242 -0.05914728716015816
storage[2822] = -13'b0000011111000; // -248 -0.060555726289749146
storage[2823] = -13'b0000110010100; // -404 -0.0985981747508049
storage[2824] =  13'b0000000011100; // 28 0.0067282491363584995
storage[2825] = -13'b0000010101011; // -171 -0.04178687185049057
storage[2826] = -13'b0000011110000; // -240 -0.05870181322097778
storage[2827] =  13'b0000011111010; // 250 0.060940586030483246
storage[2828] = -13'b0000000111010; // -58 -0.014222371391952038
storage[2829] = -13'b0000000010010; // -18 -0.004291166085749865
storage[2830] = -13'b0000000111101; // -61 -0.014907319098711014
storage[2831] =  13'b0001010101101; // 685 0.16716526448726654
storage[2832] =  13'b0001000010101; // 533 0.13001348078250885
storage[2833] = -13'b0001011001010; // -714 -0.17435233294963837
storage[2834] = -13'b0000101010101; // -341 -0.0831378772854805
storage[2835] = -13'b0000010000001; // -129 -0.031406745314598083
storage[2836] =  13'b0000010100011; // 163 0.039846476167440414
storage[2837] =  13'b0001000011110; // 542 0.13227149844169617
storage[2838] =  13'b0000111000010; // 450 0.10990579426288605
storage[2839] = -13'b0001010010001; // -657 -0.16033901274204254
storage[2840] =  13'b0000000000001; // 1 0.00016143321408890188
storage[2841] =  13'b0000001000110; // 70 0.017069265246391296
storage[2842] = -13'b0000000001101; // -13 -0.003106459276750684
storage[2843] =  13'b0000010000100; // 132 0.03211955353617668
storage[2844] =  13'b0001100010001; // 785 0.19161710143089294
storage[2845] = -13'b0000000111000; // -56 -0.013645771890878677
storage[2846] = -13'b0000001000101; // -69 -0.016827579587697983
storage[2847] = -13'b0000000011100; // -28 -0.006907626520842314
storage[2848] = -13'b0000111110000; // -496 -0.12119961529970169
storage[2849] = -13'b0000011100101; // -229 -0.055825378745794296
storage[2850] = -13'b0000010100100; // -164 -0.04010962322354317
storage[2851] =  13'b0000011000110; // 198 0.04841393232345581
storage[2852] =  13'b0000111111010; // 506 0.12358944863080978
storage[2853] = -13'b0000001001001; // -73 -0.017729666084051132
storage[2854] =  13'b0000001100010; // 98 0.023985860869288445
storage[2855] = -13'b0000101000111; // -327 -0.07992987334728241
storage[2856] =  13'b0000000100100; // 36 0.008885091170668602
storage[2857] = -13'b0010000000001; // -1025 -0.25026801228523254
storage[2858] = -13'b0001000001110; // -526 -0.12830138206481934
storage[2859] =  13'b0000101101101; // 365 0.08920362591743469
storage[2860] = -13'b0001001010111; // -599 -0.14632907509803772
storage[2861] =  13'b0000110010110; // 406 0.09920639544725418
storage[2862] =  13'b0000100100111; // 295 0.07211996614933014
storage[2863] =  13'b0001010010000; // 656 0.1601828634738922
storage[2864] =  13'b0000110010100; // 404 0.09869469702243805
storage[2865] =  13'b0000001110001; // 113 0.027487074956297874
storage[2866] = -13'b0000011101101; // -237 -0.05797076225280762
storage[2867] = -13'b0000010101110; // -174 -0.042540788650512695
storage[2868] =  13'b0000010011010; // 154 0.0375404879450798
storage[2869] = -13'b0001001111111; // -639 -0.15590707957744598
storage[2870] = -13'b0000111011010; // -474 -0.1157398596405983
storage[2871] = -13'b0000000110100; // -52 -0.012671321630477905
storage[2872] =  13'b0000001101110; // 110 0.026774032041430473
storage[2873] =  13'b0000001111010; // 122 0.029669655486941338
storage[2874] =  13'b0000001100010; // 98 0.023831570520997047
storage[2875] =  13'b0000100111110; // 318 0.0776381865143776
storage[2876] = -13'b0000000101001; // -41 -0.010093895718455315
storage[2877] = -13'b0000110110101; // -437 -0.10672944784164429
storage[2878] =  13'b0000101011111; // 351 0.08573032915592194
storage[2879] = -13'b0000001111100; // -124 -0.030316367745399475
storage[2880] =  13'b0000011000110; // 198 0.048443760722875595
storage[2881] = -13'b0000000010100; // -20 -0.004793714266270399
storage[2882] = -13'b0000000101010; // -42 -0.010247177444398403
storage[2883] = -13'b0000010101011; // -171 -0.04179145768284798
storage[2884] = -13'b0000000110001; // -49 -0.01189897209405899
storage[2885] = -13'b0000000010000; // -16 -0.0038620191626250744
storage[2886] = -13'b0000010011101; // -157 -0.038290802389383316
storage[2887] =  13'b0000010011000; // 152 0.03699495643377304
storage[2888] = -13'b0000001010111; // -87 -0.021225931122899055
storage[2889] =  13'b0000011011010; // 218 0.05333864688873291
storage[2890] = -13'b0000010101000; // -168 -0.04097599908709526
storage[2891] =  13'b0000001000100; // 68 0.016643906012177467
storage[2892] = -13'b0000001001110; // -78 -0.01910078153014183
storage[2893] = -13'b0000111000001; // -449 -0.10969598591327667
storage[2894] =  13'b0000000101011; // 43 0.010498619638383389
storage[2895] =  13'b0000100110010; // 306 0.07468477636575699
storage[2896] = -13'b0000100100000; // -288 -0.0702308788895607
storage[2897] =  13'b0000010011111; // 159 0.03872133791446686
storage[2898] =  13'b0000100010001; // 273 0.06656511127948761
storage[2899] = -13'b0000001000010; // -66 -0.016127778217196465
storage[2900] = -13'b0000001000101; // -69 -0.016875678673386574
storage[2901] =  13'b0000101101101; // 365 0.08918825536966324
storage[2902] = -13'b0000011111011; // -251 -0.061214279383420944
storage[2903] =  13'b0000101001010; // 330 0.08066299557685852
storage[2904] =  13'b0000110010000; // 400 0.09776212275028229
storage[2905] = -13'b0000110100001; // -417 -0.10177963227033615
storage[2906] =  13'b0000001001111; // 79 0.01920483633875847
storage[2907] =  13'b0000111100000; // 480 0.11728876084089279
storage[2908] =  13'b0000001000010; // 66 0.016006696969270706
storage[2909] =  13'b0000101010010; // 338 0.08241153508424759
storage[2910] =  13'b0000001000001; // 65 0.015747249126434326
storage[2911] = -13'b0000100000100; // -260 -0.06357652693986893
storage[2912] = -13'b0000100011111; // -287 -0.07006307691335678
storage[2913] =  13'b0000010110100; // 180 0.04395774379372597
storage[2914] = -13'b0000001001111; // -79 -0.019300058484077454
storage[2915] = -13'b0000010011101; // -157 -0.03823327273130417
storage[2916] =  13'b0000011000000; // 192 0.046824581921100616
storage[2917] = -13'b0000110100111; // -423 -0.1032634973526001
storage[2918] = -13'b0000111011000; // -472 -0.11527340859174728
storage[2919] = -13'b0000011000100; // -196 -0.047822173684835434
storage[2920] = -13'b0001110101100; // -940 -0.22956086695194244
storage[2921] = -13'b0001101011000; // -856 -0.20893152058124542
storage[2922] = -13'b0000011001100; // -204 -0.04982447624206543
storage[2923] = -13'b0001011011101; // -733 -0.1790146827697754
storage[2924] = -13'b0000110011110; // -414 -0.1009795144200325
storage[2925] = -13'b0000011101100; // -236 -0.057649411261081696
storage[2926] =  13'b0000000011010; // 26 0.006390304304659367
storage[2927] =  13'b0000010101111; // 175 0.042802128940820694
storage[2928] =  13'b0000001001001; // 73 0.017912795767188072
storage[2929] = -13'b0000111111001; // -505 -0.12330400198698044
storage[2930] = -13'b0000100000110; // -262 -0.06399885565042496
storage[2931] = -13'b0000101010110; // -342 -0.0836172103881836
storage[2932] = -13'b0000011000011; // -195 -0.04756933078169823
storage[2933] =  13'b0000000001010; // 10 0.0024440737906843424
storage[2934] =  13'b0000010101011; // 171 0.04168068990111351
storage[2935] =  13'b0001100100100; // 804 0.19633562862873077
storage[2936] =  13'b0000100110001; // 305 0.07444579899311066
storage[2937] = -13'b0000010000111; // -135 -0.03297464922070503
storage[2938] =  13'b0000101101101; // 365 0.08903685957193375
storage[2939] =  13'b0000110101011; // 427 0.10419680923223495
storage[2940] =  13'b0000100110110; // 310 0.07571669667959213
storage[2941] =  13'b0000010110110; // 182 0.04448087513446808
storage[2942] =  13'b0001010001110; // 654 0.15965411067008972
storage[2943] =  13'b0000011001000; // 200 0.04874521866440773
storage[2944] = -13'b0000100000011; // -259 -0.06332456320524216
storage[2945] =  13'b0000001101000; // 104 0.025345416739583015
storage[2946] =  13'b0001000100000; // 544 0.13286246359348297
storage[2947] =  13'b0000001000100; // 68 0.016528591513633728
storage[2948] =  13'b0000001010000; // 80 0.01958574913442135
storage[2949] = -13'b0000001010110; // -86 -0.020907815545797348
storage[2950] = -13'b0000011100011; // -227 -0.05533118173480034
storage[2951] = -13'b0000000010101; // -21 -0.005064947530627251
storage[2952] =  13'b0000111011000; // 472 0.11512865871191025
storage[2953] = -13'b0000011011011; // -219 -0.05357569083571434
storage[2954] =  13'b0000001011010; // 90 0.02193932980298996
storage[2955] =  13'b0000000000100; // 4 0.0010415336582809687
storage[2956] =  13'b0000011000011; // 195 0.04769274219870567
storage[2957] =  13'b0000000011000; // 24 0.005902649834752083
storage[2958] =  13'b0000011101001; // 233 0.056896913796663284
storage[2959] =  13'b0000010000000; // 128 0.03136379271745682
storage[2960] =  13'b0001000010001; // 529 0.12915991246700287
storage[2961] =  13'b0000101010101; // 341 0.08336492627859116
storage[2962] =  13'b0000010110111; // 183 0.044721074402332306
storage[2963] =  13'b0001001010011; // 595 0.1452360600233078
storage[2964] =  13'b0000100101011; // 299 0.07305930554866791
storage[2965] = -13'b0000000110010; // -50 -0.012290677055716515
storage[2966] =  13'b0000010111000; // 184 0.0448906347155571
storage[2967] =  13'b0000000000001; // 1 0.00016596396744716913
storage[2968] = -13'b0000000100100; // -36 -0.0087088318541646
storage[2969] =  13'b0000011000011; // 195 0.047574110329151154
storage[2970] =  13'b0000010011000; // 152 0.037089962512254715
storage[2971] =  13'b0000100001001; // 265 0.06465566158294678
storage[2972] =  13'b0000011011101; // 221 0.05388094112277031
storage[2973] = -13'b0000001110011; // -115 -0.028063081204891205
storage[2974] = -13'b0000101011110; // -350 -0.0853710025548935
storage[2975] =  13'b0000000100000; // 32 0.007823443971574306
storage[2976] =  13'b0000000101100; // 44 0.010782947763800621
storage[2977] = -13'b0000000100100; // -36 -0.008812964893877506
storage[2978] = -13'b0000011001011; // -203 -0.04943874105811119
storage[2979] = -13'b0000101011010; // -346 -0.08446318656206131
storage[2980] =  13'b0000100011001; // 281 0.06872440129518509
storage[2981] = -13'b0000000001001; // -9 -0.00218304805457592
storage[2982] = -13'b0000000111100; // -60 -0.014529724605381489
storage[2983] = -13'b0001000101111; // -559 -0.1363966166973114
storage[2984] = -13'b0000110010011; // -403 -0.09833361208438873
storage[2985] = -13'b0000011001110; // -206 -0.050347700715065
storage[2986] =  13'b0000110100011; // 419 0.10231778770685196
storage[2987] =  13'b0000001100100; // 100 0.024510011076927185
storage[2988] = -13'b0000000010101; // -21 -0.0050930785946547985
storage[2989] =  13'b0000010000111; // 135 0.03293134272098541
storage[2990] = -13'b0000011010110; // -214 -0.052368126809597015
storage[2991] =  13'b0000111101000; // 488 0.11903753876686096
storage[2992] = -13'b0000010101010; // -170 -0.04140021279454231
storage[2993] =  13'b0000000101100; // 44 0.010795499198138714
storage[2994] =  13'b0000001100001; // 97 0.023799054324626923
storage[2995] =  13'b0000001100110; // 102 0.024807821959257126
storage[2996] =  13'b0000011111001; // 249 0.060826510190963745
storage[2997] =  13'b0000001010100; // 84 0.020420167595148087
storage[2998] =  13'b0000000011010; // 26 0.0062893531285226345
storage[2999] = -13'b0000010101100; // -172 -0.041907381266355515
storage[3000] = -13'b0001001111101; // -637 -0.15556968748569489
storage[3001] = -13'b0000010101011; // -171 -0.04163052886724472
storage[3002] =  13'b0000001101100; // 108 0.02640056237578392
storage[3003] = -13'b0000101100010; // -354 -0.08648741990327835
storage[3004] =  13'b0000010101101; // 173 0.04225872457027435
storage[3005] =  13'b0000110000010; // 386 0.09419641643762589
storage[3006] = -13'b0000001111101; // -125 -0.030620979145169258
storage[3007] =  13'b0000010111000; // 184 0.044874198734760284
storage[3008] = -13'b0000100111101; // -317 -0.07734077423810959
storage[3009] = -13'b0000001011101; // -93 -0.02268955111503601
storage[3010] = -13'b0000001010001; // -81 -0.019878700375556946
storage[3011] =  13'b0000011100101; // 229 0.05600602924823761
storage[3012] =  13'b0000000110110; // 54 0.013172732666134834
storage[3013] =  13'b0001010100000; // 672 0.164020836353302
storage[3014] =  13'b0000110100000; // 416 0.10161468386650085
storage[3015] =  13'b0000011110001; // 241 0.058951348066329956
storage[3016] = -13'b0000010110111; // -183 -0.04457980394363403
storage[3017] = -13'b0000111110011; // -499 -0.12186450511217117
storage[3018] =  13'b0001000001000; // 520 0.12704168260097504
storage[3019] = -13'b0000101000111; // -327 -0.07984765619039536
storage[3020] = -13'b0001011000110; // -710 -0.17336063086986542
storage[3021] = -13'b0000000111101; // -61 -0.014803402125835419
storage[3022] = -13'b0000001100010; // -98 -0.024018920958042145
storage[3023] = -13'b0010011111100; // -1276 -0.3115273416042328
storage[3024] = -13'b0000011111010; // -250 -0.06096593663096428
storage[3025] = -13'b0000000101101; // -45 -0.010880823247134686
storage[3026] =  13'b0000001011011; // 91 0.02231629751622677
storage[3027] = -13'b0000001010100; // -84 -0.020582325756549835
storage[3028] = -13'b0000100100100; // -292 -0.07136428356170654
storage[3029] = -13'b0000010001001; // -137 -0.033409785479307175
storage[3030] =  13'b0000101101011; // 363 0.08868424594402313
storage[3031] = -13'b0001000010100; // -532 -0.12994620203971863
storage[3032] =  13'b0000001001010; // 74 0.017948556691408157
storage[3033] =  13'b0000100101011; // 299 0.07302025705575943
storage[3034] = -13'b0000101100110; // -358 -0.08732573688030243
storage[3035] =  13'b0000000011011; // 27 0.006629134528338909
storage[3036] = -13'b0000001101011; // -107 -0.026052795350551605
storage[3037] =  13'b0000101011010; // 346 0.08456246554851532
storage[3038] = -13'b0000000110101; // -53 -0.01282186433672905
storage[3039] = -13'b0000111000011; // -451 -0.1102244183421135
storage[3040] = -13'b0001010010011; // -659 -0.16083218157291412
storage[3041] =  13'b0000001001111; // 79 0.019370222464203835
storage[3042] =  13'b0000111110011; // 499 0.12178482115268707
storage[3043] =  13'b0000100111011; // 315 0.07693618535995483
storage[3044] = -13'b0000010110101; // -181 -0.04427868500351906
storage[3045] = -13'b0000011110010; // -242 -0.05904371663928032
storage[3046] =  13'b0000001010100; // 84 0.020507240667939186
storage[3047] = -13'b0010010010100; // -1172 -0.2861703336238861
storage[3048] = -13'b0001100111001; // -825 -0.20130085945129395
storage[3049] = -13'b0000011000000; // -192 -0.04685424268245697
storage[3050] = -13'b0001011011101; // -733 -0.1790589839220047
storage[3051] =  13'b0000011101100; // 236 0.057686977088451385
storage[3052] = -13'b0001001100111; // -615 -0.15025953948497772
storage[3053] = -13'b0000000110111; // -55 -0.01337797474116087
storage[3054] =  13'b0000101000101; // 325 0.07935018092393875
storage[3055] = -13'b0011001110010; // -1650 -0.402861624956131
storage[3056] = -13'b0000001100001; // -97 -0.023639528080821037
storage[3057] =  13'b0000011111000; // 248 0.06056418642401695
storage[3058] = -13'b0001111100001; // -993 -0.2423948049545288
storage[3059] = -13'b0000011100100; // -228 -0.05577758327126503
storage[3060] = -13'b0000000001010; // -10 -0.002419902943074703
storage[3061] = -13'b0000001000001; // -65 -0.015750553458929062
storage[3062] = -13'b0000000011100; // -28 -0.006874231155961752
storage[3063] = -13'b0000011001111; // -207 -0.050420112907886505
storage[3064] =  13'b0000010101011; // 171 0.041780948638916016
storage[3065] = -13'b0000101011010; // -346 -0.08450092375278473
storage[3066] =  13'b0000000011011; // 27 0.006626218091696501
storage[3067] = -13'b0000111111010; // -506 -0.12347038835287094
storage[3068] = -13'b0000101110111; // -375 -0.09156912565231323
storage[3069] =  13'b0000000111011; // 59 0.014483585022389889
storage[3070] =  13'b0000011111110; // 254 0.061982300132513046
storage[3071] = -13'b0000000110000; // -48 -0.011838840320706367
storage[3072] = -13'b0000011110010; // -242 -0.059078991413116455
storage[3073] =  13'b0000100001111; // 271 0.06613883376121521
storage[3074] =  13'b0000010011000; // 152 0.037127360701560974
storage[3075] = -13'b0000000001000; // -8 -0.001995360478758812
storage[3076] =  13'b0000001111011; // 123 0.030085556209087372
storage[3077] =  13'b0000010101011; // 171 0.04178180918097496
storage[3078] = -13'b0000001100010; // -98 -0.02384479157626629
storage[3079] = -13'b0000011010111; // -215 -0.05243206024169922
storage[3080] =  13'b0000000110011; // 51 0.012537401169538498
storage[3081] =  13'b0000001110000; // 112 0.02744225226342678
storage[3082] =  13'b0000011111101; // 253 0.06177873536944389
storage[3083] =  13'b0000000001110; // 14 0.0034581469371914864
storage[3084] = -13'b0000010001010; // -138 -0.03357371315360069
storage[3085] = -13'b0000000100000; // -32 -0.00772104924544692
storage[3086] = -13'b0000011101110; // -238 -0.05817796289920807
storage[3087] =  13'b0000011000101; // 197 0.048182908445596695
storage[3088] =  13'b0000010111111; // 191 0.04658155515789986
storage[3089] = -13'b0000011111000; // -248 -0.06056070327758789
storage[3090] =  13'b0000001011100; // 92 0.02248658798635006
storage[3091] = -13'b0000000110110; // -54 -0.013088797219097614
storage[3092] =  13'b0000011111011; // 251 0.061308104544878006
storage[3093] = -13'b0000100001011; // -267 -0.065268874168396
storage[3094] = -13'b0000000011100; // -28 -0.006804642733186483
storage[3095] = -13'b0000010101010; // -170 -0.04158249497413635
storage[3096] = -13'b0000101111010; // -378 -0.09227423369884491
storage[3097] =  13'b0000000000110; // 6 0.0015806981828063726
storage[3098] =  13'b0000010000110; // 134 0.03277634456753731
storage[3099] = -13'b0000101111100; // -380 -0.09282822161912918
storage[3100] = -13'b0000010010101; // -149 -0.03645223379135132
storage[3101] = -13'b0000011111001; // -249 -0.06077536195516586
storage[3102] = -13'b0010001000110; // -1094 -0.2670592963695526
storage[3103] =  13'b0000110011010; // 410 0.10014016926288605
storage[3104] =  13'b0001010011011; // 667 0.16280978918075562
storage[3105] =  13'b0000000110011; // 51 0.012406366877257824
storage[3106] =  13'b0000100010100; // 276 0.0673506036400795
storage[3107] =  13'b0000010001111; // 143 0.03498482704162598
storage[3108] = -13'b0001011111100; // -764 -0.18656659126281738
storage[3109] =  13'b0000011100111; // 231 0.05640500411391258
storage[3110] = -13'b0001010010010; // -658 -0.16060961782932281
storage[3111] = -13'b0000001111000; // -120 -0.02935878187417984
storage[3112] =  13'b0000100000100; // 260 0.06338682770729065
storage[3113] = -13'b0000001110010; // -114 -0.027822906151413918
storage[3114] =  13'b0000101001010; // 330 0.0806867703795433
storage[3115] = -13'b0000101001001; // -329 -0.08020644634962082
storage[3116] = -13'b0000011010000; // -208 -0.05070682242512703
storage[3117] = -13'b0000010110011; // -179 -0.04367451369762421
storage[3118] = -13'b0000011110111; // -247 -0.06021270900964737
storage[3119] = -13'b0000010111001; // -185 -0.04508071765303612
storage[3120] =  13'b0000010110110; // 182 0.04432094469666481
storage[3121] = -13'b0000001010000; // -80 -0.019440872594714165
storage[3122] = -13'b0000010001011; // -139 -0.03394625708460808
storage[3123] = -13'b0001010001111; // -655 -0.15999284386634827
storage[3124] = -13'b0000000101001; // -41 -0.00989177729934454
storage[3125] = -13'b0000110100010; // -418 -0.10209478437900543
storage[3126] = -13'b0000011011001; // -217 -0.05295363813638687
storage[3127] =  13'b0000010001111; // 143 0.03497328609228134
storage[3128] = -13'b0000001100011; // -99 -0.0240534208714962
storage[3129] =  13'b0000000101101; // 45 0.011104959063231945
storage[3130] =  13'b0000101100100; // 356 0.08686087280511856
storage[3131] = -13'b0000000010110; // -22 -0.005272642243653536
storage[3132] = -13'b0000100001010; // -266 -0.06482894718647003
storage[3133] = -13'b0000001101010; // -106 -0.025801856070756912
storage[3134] = -13'b0000011101111; // -239 -0.058461371809244156
storage[3135] = -13'b0000100001111; // -271 -0.06605090200901031
storage[3136] = -13'b0001101000101; // -837 -0.20435597002506256
storage[3137] = -13'b0001100001001; // -777 -0.18966129422187805
storage[3138] =  13'b0000000000100; // 4 0.0010984791442751884
storage[3139] = -13'b0000100111000; // -312 -0.07624101638793945
storage[3140] = -13'b0001001000100; // -580 -0.14158011972904205
storage[3141] = -13'b0000000110110; // -54 -0.01313759945333004
storage[3142] = -13'b0000101000110; // -326 -0.07954113930463791
storage[3143] = -13'b0000110111001; // -441 -0.1076536774635315
storage[3144] = -13'b0000010001010; // -138 -0.03371310606598854
storage[3145] = -13'b0000011101000; // -232 -0.05655533820390701
storage[3146] =  13'b0000010000100; // 132 0.03227118402719498
storage[3147] = -13'b0000000100010; // -34 -0.008284501731395721
storage[3148] =  13'b0000011100001; // 225 0.05494612827897072
storage[3149] =  13'b0000101111100; // 380 0.09268641471862793
storage[3150] = -13'b0000000011001; // -25 -0.006006804760545492
storage[3151] = -13'b0000111100010; // -482 -0.11777506023645401
storage[3152] = -13'b0000010111101; // -189 -0.046213872730731964
storage[3153] =  13'b0000011100000; // 224 0.054672155529260635
storage[3154] = -13'b0000111110001; // -497 -0.12137424200773239
storage[3155] =  13'b0000100110101; // 309 0.07535391300916672
storage[3156] =  13'b0000001000010; // 66 0.016215454787015915
storage[3157] = -13'b0000000111010; // -58 -0.014198854565620422
storage[3158] = -13'b0000101100101; // -357 -0.08719833940267563
storage[3159] = -13'b0001101110110; // -886 -0.21636469662189484
storage[3160] = -13'b0000010111011; // -187 -0.04553712159395218
storage[3161] =  13'b0000011011111; // 223 0.05445747449994087
storage[3162] = -13'b0001001100111; // -615 -0.15026657283306122
storage[3163] =  13'b0000101001011; // 331 0.080854631960392
storage[3164] =  13'b0000011011111; // 223 0.05439795181155205
storage[3165] = -13'b0000101010100; // -340 -0.08293597400188446
storage[3166] =  13'b0000110101100; // 428 0.10449245572090149
storage[3167] = -13'b0000100110010; // -306 -0.07474618405103683
storage[3168] = -13'b0000001011010; // -90 -0.02201741188764572
storage[3169] =  13'b0000111000010; // 450 0.10979996621608734
storage[3170] =  13'b0000101001100; // 332 0.08101970702409744
storage[3171] =  13'b0000000000010; // 2 0.000479805312352255
storage[3172] =  13'b0000000101011; // 43 0.010594303719699383
storage[3173] =  13'b0000100011011; // 283 0.06906396895647049
storage[3174] = -13'b0000101000101; // -325 -0.079233817756176
storage[3175] = -13'b0000000000000; // 0 -9.146129013970494e-05
storage[3176] = -13'b0000001101010; // -106 -0.025927100330591202
storage[3177] =  13'b0000001000010; // 66 0.016167987138032913
storage[3178] = -13'b0000000111001; // -57 -0.0139521025121212
storage[3179] = -13'b0000001011011; // -91 -0.02220519818365574
storage[3180] = -13'b0000101110110; // -374 -0.09141910821199417
storage[3181] =  13'b0000111110011; // 499 0.1217595711350441
storage[3182] = -13'b0000000010111; // -23 -0.005515394266694784
storage[3183] =  13'b0000101100000; // 352 0.0858457013964653
storage[3184] =  13'b0000101101110; // 366 0.08939771354198456
storage[3185] = -13'b0010111101010; // -1514 -0.3697243630886078
storage[3186] =  13'b0001111101111; // 1007 0.24583926796913147
storage[3187] =  13'b0000010111010; // 186 0.045328784734010696
storage[3188] =  13'b0000010011101; // 157 0.03822833672165871
storage[3189] = -13'b0000001010010; // -82 -0.020052464678883553
storage[3190] =  13'b0000011110100; // 244 0.05959874019026756
storage[3191] =  13'b0000001000010; // 66 0.016126492992043495
storage[3192] =  13'b0000011100101; // 229 0.05594636872410774
storage[3193] = -13'b0001000111110; // -574 -0.14006228744983673
storage[3194] = -13'b0000111000101; // -453 -0.11058869957923889
storage[3195] = -13'b0001000010110; // -534 -0.13031375408172607
storage[3196] = -13'b0000000010110; // -22 -0.005362862255424261
storage[3197] =  13'b0000011001001; // 201 0.049178287386894226
storage[3198] =  13'b0000011100110; // 230 0.056267280131578445
storage[3199] = -13'b0000000110100; // -52 -0.012637716718018055
storage[3200] = -13'b0011101110101; // -1909 -0.46599870920181274
storage[3201] = -13'b0000111111001; // -505 -0.12320943921804428
storage[3202] =  13'b0000011110110; // 246 0.06014710292220116
storage[3203] = -13'b0010100110101; // -1333 -0.325454443693161
storage[3204] =  13'b0001111001011; // 971 0.23698410391807556
storage[3205] =  13'b0000100100010; // 290 0.07068856805562973
storage[3206] =  13'b0000100000110; // 262 0.0639519914984703
storage[3207] =  13'b0000001101100; // 108 0.026476241648197174
storage[3208] =  13'b0000001001101; // 77 0.018874336034059525
storage[3209] = -13'b0000000011000; // -24 -0.005798249505460262
storage[3210] = -13'b0000011011101; // -221 -0.05393649637699127
storage[3211] = -13'b0000000010101; // -21 -0.005194821860641241
storage[3212] =  13'b0000001110011; // 115 0.028175514191389084
storage[3213] = -13'b0000011111000; // -248 -0.06046596169471741
storage[3214] = -13'b0000000010110; // -22 -0.005488619673997164
storage[3215] =  13'b0000000011000; // 24 0.005788235459476709
storage[3216] =  13'b0000101010100; // 340 0.08307871222496033
storage[3217] = -13'b0000100011110; // -286 -0.06987232714891434
storage[3218] =  13'b0000101010000; // 336 0.08194270730018616
storage[3219] =  13'b0000110000011; // 387 0.09456528723239899
storage[3220] = -13'b0001000010100; // -532 -0.12998038530349731
storage[3221] = -13'b0000000111001; // -57 -0.013927157036960125
storage[3222] =  13'b0000110010101; // 405 0.09891210496425629
storage[3223] = -13'b0000010110110; // -182 -0.044311754405498505
storage[3224] = -13'b0000001000100; // -68 -0.01669529266655445
storage[3225] =  13'b0000101000111; // 327 0.07971882075071335
storage[3226] =  13'b0000001011100; // 92 0.02253318764269352
storage[3227] =  13'b0000001010011; // 83 0.020152952522039413
storage[3228] =  13'b0000001010110; // 86 0.02096700295805931
storage[3229] =  13'b0000001001101; // 77 0.018751021474599838
storage[3230] =  13'b0000000010000; // 16 0.004007733892649412
storage[3231] = -13'b0000100001100; // -268 -0.06542510539293289
storage[3232] = -13'b0000011001110; // -206 -0.05026150122284889
storage[3233] =  13'b0000000011101; // 29 0.007099532522261143
storage[3234] =  13'b0000001010011; // 83 0.020299995318055153
storage[3235] = -13'b0000110011111; // -415 -0.10138186067342758
storage[3236] = -13'b0000000011101; // -29 -0.00716381287202239
storage[3237] =  13'b0000010110001; // 177 0.043103061616420746
storage[3238] = -13'b0001110100000; // -928 -0.22657974064350128
storage[3239] = -13'b0000010101110; // -174 -0.04237636178731918
storage[3240] = -13'b0000101011010; // -346 -0.08440161496400833
storage[3241] =  13'b0000000011000; // 24 0.005819160025566816
storage[3242] =  13'b0000100011011; // 283 0.06913884729146957
storage[3243] =  13'b0000000110101; // 53 0.012972152791917324
storage[3244] = -13'b0000000001000; // -8 -0.0020606648176908493
storage[3245] = -13'b0000010111000; // -184 -0.0448710173368454
storage[3246] =  13'b0000110101000; // 424 0.10357403010129929
storage[3247] = -13'b0000010111011; // -187 -0.04553527384996414
storage[3248] = -13'b0000001100011; // -99 -0.024148231372237206
storage[3249] =  13'b0000010001101; // 141 0.034421682357788086
storage[3250] = -13'b0000000100011; // -35 -0.008477800525724888
storage[3251] =  13'b0000001001101; // 77 0.01879037544131279
storage[3252] =  13'b0000001001101; // 77 0.018880443647503853
storage[3253] = -13'b0000011111111; // -255 -0.06224583461880684
storage[3254] = -13'b0000011100111; // -231 -0.05632294714450836
storage[3255] = -13'b0001010110010; // -690 -0.16848541796207428
storage[3256] =  13'b0000000001111; // 15 0.00369332660920918
storage[3257] = -13'b0000100101111; // -303 -0.07387075573205948
storage[3258] = -13'b0000111000100; // -452 -0.1102437898516655
storage[3259] = -13'b0000000101110; // -46 -0.011313263326883316
storage[3260] = -13'b0000100100101; // -293 -0.07161016762256622
storage[3261] = -13'b0001010111000; // -696 -0.16993629932403564
storage[3262] =  13'b0000000011010; // 26 0.006261416245251894
storage[3263] = -13'b0000111001100; // -460 -0.11223427206277847
storage[3264] = -13'b0000011110001; // -241 -0.058901943266391754
storage[3265] =  13'b0000001111100; // 124 0.030332209542393684
storage[3266] =  13'b0000011011001; // 217 0.05291195213794708
storage[3267] =  13'b0000011001110; // 206 0.05026834458112717
storage[3268] = -13'b0000111000001; // -449 -0.10956012457609177
storage[3269] =  13'b0000010110000; // 176 0.042964208871126175
storage[3270] = -13'b0000000110001; // -49 -0.011846532113850117
storage[3271] =  13'b0000011110101; // 245 0.059890132397413254
storage[3272] = -13'b0001000001010; // -522 -0.1273622214794159
storage[3273] = -13'b0001000110000; // -560 -0.13677595555782318
storage[3274] = -13'b0000100001110; // -270 -0.06586244702339172
storage[3275] = -13'b0000100111011; // -315 -0.07683029770851135
storage[3276] =  13'b0000001011010; // 90 0.021991858258843422
storage[3277] =  13'b0000110000011; // 387 0.09448004513978958
storage[3278] = -13'b0000010011001; // -153 -0.0373050831258297
storage[3279] = -13'b0000001010110; // -86 -0.020903419703245163
storage[3280] =  13'b0000010000010; // 130 0.031675584614276886
storage[3281] =  13'b0000010101011; // 171 0.04168105497956276
storage[3282] =  13'b0000001100001; // 97 0.023723537102341652
storage[3283] = -13'b0000101110101; // -373 -0.0911017581820488
storage[3284] = -13'b0000000000100; // -4 -0.0009406586177647114
storage[3285] =  13'b0000010111011; // 187 0.04565434530377388
storage[3286] =  13'b0001000001110; // 526 0.12850691378116608
storage[3287] =  13'b0000101100101; // 357 0.08716394752264023
storage[3288] =  13'b0000001011111; // 95 0.02307247556746006
storage[3289] = -13'b0001000011010; // -538 -0.13124389946460724
storage[3290] = -13'b0000101000100; // -324 -0.07900644838809967
storage[3291] =  13'b0000001100011; // 99 0.024117687717080116
storage[3292] = -13'b0000011100011; // -227 -0.05536244064569473
storage[3293] = -13'b0000010111101; // -189 -0.046027787029743195
storage[3294] =  13'b0000011101110; // 238 0.05817323923110962
storage[3295] =  13'b0000101110111; // 375 0.0915687307715416
storage[3296] = -13'b0000100010101; // -277 -0.06770350784063339
storage[3297] = -13'b0000100100000; // -288 -0.0702924057841301
storage[3298] = -13'b0000110001011; // -395 -0.09644988924264908
storage[3299] = -13'b0000011011011; // -219 -0.05336529761552811
storage[3300] =  13'b0000010110000; // 176 0.0430198535323143
storage[3301] =  13'b0000000000011; // 3 0.0008130369824357331
storage[3302] =  13'b0000001001111; // 79 0.019367871806025505
storage[3303] =  13'b0000100010101; // 277 0.06765076518058777
storage[3304] = -13'b0000101001101; // -333 -0.08135708421468735
storage[3305] = -13'b0000000100111; // -39 -0.009501686319708824
storage[3306] =  13'b0000100111111; // 319 0.07783612608909607
storage[3307] =  13'b0000100010101; // 277 0.06751368939876556
storage[3308] =  13'b0000000011010; // 26 0.006289046257734299
storage[3309] =  13'b0000001000110; // 70 0.017025543376803398
storage[3310] =  13'b0000111011011; // 475 0.11587739735841751
storage[3311] =  13'b0000001011001; // 89 0.021777847781777382
storage[3312] = -13'b0001001010110; // -598 -0.1459764689207077
storage[3313] = -13'b0000100111110; // -318 -0.07756514102220535
storage[3314] = -13'b0000000110100; // -52 -0.012593904510140419
storage[3315] =  13'b0000001110000; // 112 0.02745850197970867
storage[3316] =  13'b0000100110111; // 311 0.07588417828083038
storage[3317] =  13'b0000100111111; // 319 0.07791142910718918
storage[3318] =  13'b0000110111101; // 445 0.10864460468292236
storage[3319] =  13'b0000100001000; // 264 0.06437386572360992
storage[3320] = -13'b0000000011101; // -29 -0.007142219226807356
storage[3321] = -13'b0000000010010; // -18 -0.004352628719061613
storage[3322] = -13'b0000011001011; // -203 -0.04945668578147888
storage[3323] = -13'b0000100000000; // -256 -0.06239677593111992
storage[3324] = -13'b0000001101011; // -107 -0.02602733112871647
storage[3325] = -13'b0001010011101; // -669 -0.16321739554405212
storage[3326] = -13'b0000110010010; // -402 -0.09805223345756531
storage[3327] = -13'b0000011011111; // -223 -0.05436243116855621
storage[3328] =  13'b0000001110110; // 118 0.028820456936955452
storage[3329] = -13'b0000010100010; // -162 -0.03964828699827194
storage[3330] =  13'b0000001010101; // 85 0.020665651187300682
storage[3331] =  13'b0000000101000; // 40 0.009666220284998417
storage[3332] =  13'b0000000001100; // 12 0.0029285000637173653
storage[3333] =  13'b0000011000001; // 193 0.04718094691634178
storage[3334] =  13'b0000000000011; // 3 0.000701840384863317
storage[3335] =  13'b0000001011110; // 94 0.023038992658257484
storage[3336] =  13'b0000000101100; // 44 0.010816950350999832
storage[3337] =  13'b0001000101010; // 554 0.13532941043376923
storage[3338] = -13'b0000001000000; // -64 -0.015542063862085342
storage[3339] = -13'b0000010001010; // -138 -0.03380236402153969
storage[3340] = -13'b0001000010000; // -528 -0.12893569469451904
storage[3341] = -13'b0000001000000; // -64 -0.01574467122554779
storage[3342] = -13'b0001001111011; // -635 -0.15514761209487915
storage[3343] = -13'b0000000100000; // -32 -0.007736430503427982
storage[3344] =  13'b0000101110110; // 374 0.09134361147880554
storage[3345] =  13'b0000100001110; // 270 0.06586696952581406
storage[3346] = -13'b0000010010100; // -148 -0.03603541851043701
storage[3347] = -13'b0000101000101; // -325 -0.0794065073132515
storage[3348] = -13'b0001011111001; // -761 -0.18581241369247437
storage[3349] = -13'b0000111100001; // -481 -0.11743544787168503
storage[3350] = -13'b0000000001101; // -13 -0.0031374581158161163
storage[3351] =  13'b0000100011010; // 282 0.06893635541200638
storage[3352] =  13'b0000100100010; // 290 0.07088703662157059
storage[3353] =  13'b0000110101110; // 430 0.10495816171169281
storage[3354] =  13'b0000110110000; // 432 0.10539881139993668
storage[3355] =  13'b0000010101101; // 173 0.04217527434229851
storage[3356] =  13'b0000001010010; // 82 0.02000615745782852
storage[3357] =  13'b0000100000100; // 260 0.06352292746305466
storage[3358] =  13'b0000110101001; // 425 0.10372406989336014
storage[3359] =  13'b0000100000100; // 260 0.06351085007190704
storage[3360] =  13'b0000001110001; // 113 0.027698004618287086
storage[3361] = -13'b0000010100111; // -167 -0.04069070145487785
storage[3362] = -13'b0000011100001; // -225 -0.054865676909685135
storage[3363] =  13'b0000011000010; // 194 0.047473661601543427
storage[3364] =  13'b0000011001110; // 206 0.050278641283512115
storage[3365] =  13'b0000100011010; // 282 0.06886285543441772
storage[3366] =  13'b0000011000011; // 195 0.047709837555885315
storage[3367] =  13'b0000000000110; // 6 0.0013778425054624677
storage[3368] =  13'b0000001010111; // 87 0.021279020234942436
storage[3369] = -13'b0000100110101; // -309 -0.07555316388607025
storage[3370] =  13'b0000000110101; // 53 0.013047597371041775
storage[3371] = -13'b0000001001100; // -76 -0.018478350713849068
storage[3372] = -13'b0000001110011; // -115 -0.027989698573946953
storage[3373] =  13'b0000001011011; // 91 0.02214926667511463
storage[3374] = -13'b0001000011110; // -542 -0.13235189020633698
storage[3375] = -13'b0000011000011; // -195 -0.047571346163749695
storage[3376] = -13'b0000000011010; // -26 -0.006391284521669149
storage[3377] =  13'b0000001011100; // 92 0.02249489538371563
storage[3378] =  13'b0000101111011; // 379 0.09247951954603195
storage[3379] = -13'b0000101100010; // -354 -0.08651670813560486
storage[3380] =  13'b0000000101011; // 43 0.010588839650154114
storage[3381] =  13'b0000000001001; // 9 0.002108874963596463
storage[3382] =  13'b0000010111110; // 190 0.04630151391029358
storage[3383] =  13'b0000101001110; // 334 0.08143578469753265
storage[3384] =  13'b0000101001000; // 328 0.08013346046209335
storage[3385] = -13'b0000011001011; // -203 -0.04955268278717995
storage[3386] = -13'b0000000010011; // -19 -0.0045975069515407085
storage[3387] = -13'b0000001100000; // -96 -0.023323265835642815
storage[3388] =  13'b0000101101110; // 366 0.08927187323570251
storage[3389] =  13'b0000000011101; // 29 0.007089280057698488
storage[3390] = -13'b0000010001110; // -142 -0.03464049473404884
storage[3391] = -13'b0000000010110; // -22 -0.005281451158225536
storage[3392] =  13'b0000000101010; // 42 0.010313826613128185
storage[3393] =  13'b0000011100110; // 230 0.056064214557409286
storage[3394] =  13'b0000001010110; // 86 0.021084971725940704
storage[3395] = -13'b0000000010010; // -18 -0.004339416045695543
storage[3396] = -13'b0000001011001; // -89 -0.021766113117337227
storage[3397] =  13'b0000110101011; // 427 0.10430419445037842
storage[3398] =  13'b0000101110001; // 369 0.08996766805648804
storage[3399] =  13'b0000001000111; // 71 0.017366334795951843
storage[3400] = -13'b0000001111000; // -120 -0.029200777411460876
storage[3401] = -13'b0000010001010; // -138 -0.03363335505127907
storage[3402] = -13'b0000110101110; // -430 -0.10503125190734863
storage[3403] =  13'b0000001111111; // 127 0.030949657782912254
storage[3404] =  13'b0000011010101; // 213 0.051890578120946884
storage[3405] = -13'b0000100001100; // -268 -0.06552868336439133
storage[3406] = -13'b0000011000110; // -198 -0.04839044064283371
storage[3407] = -13'b0000011010110; // -214 -0.05218829959630966
storage[3408] =  13'b0000000101101; // 45 0.010942980647087097
storage[3409] = -13'b0000100110111; // -311 -0.07591994106769562
storage[3410] =  13'b0000001000011; // 67 0.01636625826358795
storage[3411] = -13'b0000100110010; // -306 -0.07464674860239029
storage[3412] = -13'b0000010110011; // -179 -0.043699897825717926
storage[3413] = -13'b0001100000000; // -768 -0.18744227290153503
storage[3414] =  13'b0000100011010; // 282 0.06895436346530914
storage[3415] = -13'b0000001001110; // -78 -0.018924323841929436
storage[3416] = -13'b0000010100110; // -166 -0.04040973633527756
storage[3417] = -13'b0000001100111; // -103 -0.02508797124028206
storage[3418] = -13'b0001010111110; // -702 -0.17137925326824188
storage[3419] = -13'b0001001000110; // -582 -0.14199188351631165
storage[3420] = -13'b0000010010111; // -151 -0.03679807484149933
storage[3421] = -13'b0000011011011; // -219 -0.05354800820350647
storage[3422] = -13'b0000010100000; // -160 -0.039100468158721924
storage[3423] = -13'b0000011010101; // -213 -0.051893964409828186
storage[3424] =  13'b0000000110111; // 55 0.013306514360010624
storage[3425] =  13'b0000001011101; // 93 0.022605912759900093
storage[3426] =  13'b0000101111001; // 377 0.09215965121984482
storage[3427] =  13'b0000010100100; // 164 0.04007213935256004
storage[3428] =  13'b0000001111011; // 123 0.029936853796243668
storage[3429] =  13'b0000000001011; // 11 0.0025720414705574512
storage[3430] = -13'b0000000010000; // -16 -0.003902381518855691
storage[3431] =  13'b0000101011000; // 344 0.08398666232824326
storage[3432] =  13'b0000100101010; // 298 0.0728600025177002
storage[3433] =  13'b0000001100101; // 101 0.024567486718297005
storage[3434] =  13'b0000101110011; // 371 0.0905052199959755
storage[3435] =  13'b0000000011000; // 24 0.0059660556726157665
storage[3436] = -13'b0000110000000; // -384 -0.0936291366815567
storage[3437] = -13'b0001001110010; // -626 -0.15284617245197296
storage[3438] = -13'b0000000011111; // -31 -0.007520134560763836
storage[3439] =  13'b0000000100110; // 38 0.009381922893226147
storage[3440] = -13'b0000001001101; // -77 -0.01881633885204792
storage[3441] = -13'b0001000010101; // -533 -0.13013707101345062
storage[3442] =  13'b0000110001000; // 392 0.0956939160823822
storage[3443] = -13'b0001101110111; // -887 -0.21655869483947754
storage[3444] = -13'b0001010110001; // -689 -0.16831061244010925
storage[3445] =  13'b0000110111101; // 445 0.10864224284887314
storage[3446] = -13'b0000001110001; // -113 -0.027537500485777855
storage[3447] =  13'b0000100001010; // 266 0.06485992670059204
storage[3448] =  13'b0000010110101; // 181 0.044271960854530334
storage[3449] = -13'b0000111110111; // -503 -0.12269466370344162
storage[3450] = -13'b0001000100001; // -545 -0.13294488191604614
storage[3451] = -13'b0000001000110; // -70 -0.017170768231153488
storage[3452] =  13'b0000000001000; // 8 0.001967773539945483
storage[3453] = -13'b0000011101001; // -233 -0.05683257058262825
storage[3454] =  13'b0000011011110; // 222 0.054122164845466614
storage[3455] =  13'b0001101001010; // 842 0.20562151074409485
storage[3456] =  13'b0000111011110; // 478 0.11658890545368195
storage[3457] =  13'b0000100100011; // 291 0.07100847363471985
storage[3458] = -13'b0000001000001; // -65 -0.015866681933403015
storage[3459] =  13'b0000100010100; // 276 0.067457415163517
storage[3460] = -13'b0000010010101; // -149 -0.03641420602798462
storage[3461] = -13'b0000011110100; // -244 -0.05945034697651863
storage[3462] =  13'b0000101100001; // 353 0.08615602552890778
storage[3463] = -13'b0000001111010; // -122 -0.029896719381213188
storage[3464] = -13'b0001110011010; // -922 -0.22502945363521576
storage[3465] = -13'b0001100110000; // -816 -0.19920285046100616
storage[3466] =  13'b0000110010110; // 406 0.09921390563249588
storage[3467] = -13'b0000010011011; // -155 -0.037799011915922165
storage[3468] =  13'b0000011101110; // 238 0.058117639273405075
storage[3469] = -13'b0000111110000; // -496 -0.12115936726331711
storage[3470] = -13'b0001100001101; // -781 -0.190669447183609
storage[3471] = -13'b0000000110000; // -48 -0.01164384838193655
storage[3472] = -13'b0000000000100; // -4 -0.0009666372206993401
storage[3473] =  13'b0000000100001; // 33 0.007975113578140736
storage[3474] = -13'b0000010111101; // -189 -0.046138569712638855
storage[3475] =  13'b0000010000110; // 134 0.03269846364855766
storage[3476] =  13'b0000001001111; // 79 0.019363783299922943
storage[3477] =  13'b0000000000101; // 5 0.0012525392230600119
storage[3478] = -13'b0000100100001; // -289 -0.0706786960363388
storage[3479] =  13'b0000010101000; // 168 0.04107197746634483
storage[3480] =  13'b0000001110110; // 118 0.02879069186747074
storage[3481] = -13'b0000100101111; // -303 -0.07398606091737747
storage[3482] = -13'b0000010110010; // -178 -0.0434165857732296
storage[3483] = -13'b0000000110000; // -48 -0.011734604835510254
storage[3484] = -13'b0000001000110; // -70 -0.01711842603981495
storage[3485] = -13'b0001000111110; // -574 -0.14015468955039978
storage[3486] = -13'b0000010101110; // -174 -0.0424995981156826
storage[3487] =  13'b0000000101111; // 47 0.011385603807866573
storage[3488] = -13'b0000001101100; // -108 -0.026367152109742165
storage[3489] = -13'b0000001010110; // -86 -0.021031316369771957
storage[3490] =  13'b0000000010011; // 19 0.00464408565312624
storage[3491] = -13'b0001000111110; // -574 -0.1402088850736618
storage[3492] = -13'b0001010001110; // -654 -0.15955136716365814
storage[3493] = -13'b0000110011101; // -413 -0.10094653069972992
storage[3494] = -13'b0000001000010; // -66 -0.01606537215411663
storage[3495] =  13'b0000000111110; // 62 0.015020322054624557
storage[3496] = -13'b0000010000111; // -135 -0.03303862363100052
storage[3497] =  13'b0000001001101; // 77 0.01878509111702442
storage[3498] =  13'b0000010001010; // 138 0.033764198422431946
storage[3499] =  13'b0000100100101; // 293 0.07150264829397202
storage[3500] =  13'b0000000001001; // 9 0.0022488704416900873
storage[3501] = -13'b0000000010110; // -22 -0.005484444554895163
storage[3502] = -13'b0000001010000; // -80 -0.019562477245926857
storage[3503] =  13'b0000110100111; // 423 0.10336251556873322
storage[3504] =  13'b0000001100111; // 103 0.025051355361938477
storage[3505] =  13'b0000001101010; // 106 0.02583688497543335
storage[3506] =  13'b0000100101000; // 296 0.07228372991085052
storage[3507] =  13'b0000001101100; // 108 0.02633158676326275
storage[3508] =  13'b0000000110011; // 51 0.01248125359416008
storage[3509] =  13'b0000011101000; // 232 0.056756392121315
storage[3510] = -13'b0000001101111; // -111 -0.02718624845147133
storage[3511] =  13'b0000010010011; // 147 0.03595094755291939
storage[3512] =  13'b0000001000110; // 70 0.017085783183574677
storage[3513] = -13'b0001110001100; // -908 -0.22171762585639954
storage[3514] =  13'b0000000001001; // 9 0.002275089267641306
storage[3515] = -13'b0000001001110; // -78 -0.019163021817803383
storage[3516] =  13'b0000010001110; // 142 0.03469749540090561
storage[3517] =  13'b0000010011001; // 153 0.037377092987298965
storage[3518] =  13'b0000001110011; // 115 0.028119314461946487
storage[3519] =  13'b0000100100001; // 289 0.07063502073287964
storage[3520] =  13'b0000011010001; // 209 0.05103989690542221
storage[3521] =  13'b0000100101001; // 297 0.07255889475345612
storage[3522] =  13'b0000000001100; // 12 0.003050935920327902
storage[3523] = -13'b0000001101110; // -110 -0.026841912418603897
storage[3524] =  13'b0000001000101; // 69 0.016761088743805885
storage[3525] = -13'b0000101001100; // -332 -0.08105643093585968
storage[3526] = -13'b0000101101110; // -366 -0.08936721831560135
storage[3527] =  13'b0000010101111; // 175 0.042785532772541046
storage[3528] =  13'b0000111010110; // 470 0.11482195556163788
storage[3529] = -13'b0000011100100; // -228 -0.055723223835229874
storage[3530] = -13'b0000110111001; // -441 -0.1077650636434555
storage[3531] = -13'b0000010001110; // -142 -0.03465097397565842
storage[3532] =  13'b0000001111100; // 124 0.03020760416984558
storage[3533] = -13'b0000000100000; // -32 -0.007702532224357128
storage[3534] = -13'b0000000010111; // -23 -0.005715617444366217
storage[3535] =  13'b0001101011010; // 858 0.20940090715885162
storage[3536] =  13'b0001000011000; // 536 0.1308344006538391
storage[3537] =  13'b0000101011001; // 345 0.08424478769302368
storage[3538] = -13'b0000100001100; // -268 -0.06539551913738251
storage[3539] = -13'b0000100101101; // -301 -0.07341038435697556
storage[3540] =  13'b0000000001111; // 15 0.0035701037850230932
storage[3541] =  13'b0001000000011; // 515 0.1257072538137436
storage[3542] =  13'b0000001111111; // 127 0.03092244453728199
storage[3543] =  13'b0000101111001; // 377 0.09199479222297668
storage[3544] =  13'b0000000101010; // 42 0.010189519263803959
storage[3545] = -13'b0000001110100; // -116 -0.028426826000213623
storage[3546] = -13'b0000000001110; // -14 -0.003525253850966692
storage[3547] =  13'b0000000001011; // 11 0.0026817985344678164
storage[3548] = -13'b0000001000011; // -67 -0.016367604956030846
storage[3549] = -13'b0000000111001; // -57 -0.013864891603589058
storage[3550] = -13'b0000000101010; // -42 -0.010198518633842468
storage[3551] =  13'b0000001101001; // 105 0.02554984577000141
storage[3552] =  13'b0000011110000; // 240 0.0585663877427578
storage[3553] = -13'b0000110101101; // -429 -0.1047266498208046
storage[3554] = -13'b0000110001010; // -394 -0.09613484144210815
storage[3555] = -13'b0000000110110; // -54 -0.013271377421915531
storage[3556] = -13'b0000010000111; // -135 -0.03289078548550606
storage[3557] = -13'b0001000001100; // -524 -0.1279902309179306
storage[3558] = -13'b0000001111011; // -123 -0.029991626739501953
storage[3559] = -13'b0000101001100; // -332 -0.08105010539293289
storage[3560] = -13'b0001100010110; // -790 -0.1927950531244278
storage[3561] = -13'b0001000111101; // -573 -0.14000438153743744
storage[3562] = -13'b0001111010111; // -983 -0.23999442160129547
storage[3563] = -13'b0010000111101; // -1085 -0.26486480236053467
storage[3564] = -13'b0000101000010; // -322 -0.0785142108798027
storage[3565] =  13'b0000011001100; // 204 0.049800772219896317
storage[3566] =  13'b0000010101110; // 174 0.04244508966803551
storage[3567] =  13'b0000001001010; // 74 0.018177170306444168
storage[3568] = -13'b0000100110100; // -308 -0.075100839138031
storage[3569] = -13'b0000000001101; // -13 -0.0031388490460813046
storage[3570] =  13'b0000011101000; // 232 0.056724242866039276
storage[3571] = -13'b0000010010101; // -149 -0.0362984873354435
storage[3572] = -13'b0000010100100; // -164 -0.04001810401678085
storage[3573] =  13'b0000101011011; // 347 0.08471174538135529
storage[3574] = -13'b0001001101110; // -622 -0.15175266563892365
storage[3575] = -13'b0001000000111; // -519 -0.12680929899215698
storage[3576] =  13'b0000001101100; // 108 0.026318540796637535
storage[3577] = -13'b0000010000000; // -128 -0.031334083527326584
storage[3578] =  13'b0000000101011; // 43 0.010426938533782959
storage[3579] =  13'b0000100111111; // 319 0.07798943668603897
storage[3580] =  13'b0000011010010; // 210 0.051270533353090286
storage[3581] =  13'b0000001111100; // 124 0.030391262844204903
storage[3582] = -13'b0000100101000; // -296 -0.0721663311123848
storage[3583] = -13'b0001000001000; // -520 -0.12701138854026794
storage[3584] =  13'b0000010010000; // 144 0.035120848566293716
storage[3585] = -13'b0000011111000; // -248 -0.060557011514902115
storage[3586] = -13'b0001101001101; // -845 -0.20639197528362274
storage[3587] = -13'b0001010100111; // -679 -0.16579575836658478
storage[3588] = -13'b0000010110011; // -179 -0.04373258352279663
storage[3589] = -13'b0000000101011; // -43 -0.010476004332304
storage[3590] =  13'b0000100101111; // 303 0.07390716671943665
storage[3591] =  13'b0000100000001; // 257 0.06270021945238113
storage[3592] = -13'b0000101111010; // -378 -0.09230145812034607
storage[3593] = -13'b0001001011010; // -602 -0.1468837559223175
storage[3594] = -13'b0000110111001; // -441 -0.10760009288787842
storage[3595] =  13'b0000100100001; // 289 0.07060360908508301
storage[3596] =  13'b0000110011100; // 412 0.10049600154161453
storage[3597] = -13'b0001001111110; // -638 -0.15588121116161346
storage[3598] = -13'b0000001111111; // -127 -0.03095792979001999
storage[3599] =  13'b0000000001110; // 14 0.0034722741693258286
storage[3600] =  13'b0000011000010; // 194 0.047419480979442596
storage[3601] = -13'b0000100010111; // -279 -0.06816656142473221
storage[3602] = -13'b0000000000101; // -5 -0.001277462113648653
storage[3603] = -13'b0000001011101; // -93 -0.022684214636683464
storage[3604] =  13'b0000000111001; // 57 0.013872670009732246
storage[3605] = -13'b0000000011100; // -28 -0.0068896012380719185
storage[3606] =  13'b0000010001011; // 139 0.034057166427373886
storage[3607] = -13'b0000000110110; // -54 -0.013155132532119751
storage[3608] = -13'b0000011110100; // -244 -0.059475213289260864
storage[3609] = -13'b0000111010100; // -468 -0.11437363922595978
storage[3610] =  13'b0000001101001; // 105 0.02566353604197502
storage[3611] = -13'b0000001100000; // -96 -0.023316286504268646
storage[3612] = -13'b0000011011100; // -220 -0.05379675701260567
storage[3613] = -13'b0000000100110; // -38 -0.009190838783979416
storage[3614] = -13'b0000010001100; // -140 -0.03423931077122688
storage[3615] =  13'b0000001011010; // 90 0.022006770595908165
storage[3616] =  13'b0000100101000; // 296 0.07220999896526337
storage[3617] = -13'b0000000110001; // -49 -0.012041432783007622
storage[3618] =  13'b0000011110010; // 242 0.05896688625216484
storage[3619] =  13'b0000101110100; // 372 0.09094182401895523
storage[3620] =  13'b0000011101011; // 235 0.05737605318427086
storage[3621] = -13'b0001001000000; // -576 -0.14056703448295593
storage[3622] =  13'b0000010101011; // 171 0.041655246168375015
storage[3623] =  13'b0000001101100; // 108 0.026402419432997704
storage[3624] =  13'b0000000111101; // 61 0.014787392690777779
storage[3625] = -13'b0000000000001; // -1 -0.0003140512853860855
storage[3626] =  13'b0000010010101; // 149 0.03636237606406212
storage[3627] =  13'b0000000111111; // 63 0.015416346490383148
storage[3628] =  13'b0000001001100; // 76 0.018641185015439987
storage[3629] =  13'b0000000010010; // 18 0.004429843742400408
storage[3630] =  13'b0000101010011; // 339 0.08268263936042786
storage[3631] =  13'b0000100000001; // 257 0.06283356994390488
storage[3632] = -13'b0000001111100; // -124 -0.03016400709748268
storage[3633] =  13'b0000010110011; // 179 0.043639857321977615
storage[3634] =  13'b0000001010011; // 83 0.020273156464099884
storage[3635] = -13'b0001000111111; // -575 -0.14034265279769897
storage[3636] = -13'b0000100100011; // -291 -0.07105795294046402
storage[3637] = -13'b0000101011001; // -345 -0.08415667712688446
storage[3638] = -13'b0000000111110; // -62 -0.015130143612623215
storage[3639] =  13'b0000011010100; // 212 0.05184312164783478
storage[3640] =  13'b0000010100001; // 161 0.039354339241981506
storage[3641] =  13'b0000110001001; // 393 0.09595555067062378
storage[3642] =  13'b0000110111101; // 445 0.10863932222127914
storage[3643] = -13'b0000001001000; // -72 -0.017650684341788292
storage[3644] =  13'b0000001010001; // 81 0.019710645079612732
storage[3645] = -13'b0000100000100; // -260 -0.06354133784770966
storage[3646] = -13'b0000011111001; // -249 -0.06070845201611519
storage[3647] = -13'b0001001011100; // -604 -0.14741984009742737
storage[3648] = -13'b0010011000110; // -1222 -0.298279345035553
storage[3649] = -13'b0000010000110; // -134 -0.0328313410282135
storage[3650] =  13'b0000100111101; // 317 0.07736331969499588
storage[3651] =  13'b0000010100101; // 165 0.040321070700883865
storage[3652] =  13'b0000010101101; // 173 0.04220540449023247
storage[3653] =  13'b0001000001110; // 526 0.12837901711463928
storage[3654] =  13'b0000000110100; // 52 0.012798380106687546
storage[3655] = -13'b0000001101011; // -107 -0.02604791894555092
storage[3656] =  13'b0000000110110; // 54 0.013178158551454544
storage[3657] = -13'b0000101011001; // -345 -0.08434431254863739
storage[3658] =  13'b0000111101111; // 495 0.1207355484366417
storage[3659] =  13'b0000110011001; // 409 0.09986874461174011
storage[3660] = -13'b0000000110101; // -53 -0.012960975989699364
storage[3661] =  13'b0000000011000; // 24 0.005941626150161028
storage[3662] =  13'b0001010111010; // 698 0.17037507891654968
storage[3663] =  13'b0001001100111; // 615 0.1500968337059021
storage[3664] = -13'b0000100000010; // -258 -0.0629580095410347
storage[3665] = -13'b0000001010111; // -87 -0.02127683162689209
storage[3666] =  13'b0000010110001; // 177 0.04312380775809288
storage[3667] = -13'b0000010101010; // -170 -0.04149872809648514
storage[3668] =  13'b0000010011010; // 154 0.03763397037982941
storage[3669] =  13'b0000000000101; // 5 0.0013370749074965715
storage[3670] =  13'b0000001111110; // 126 0.030769772827625275
storage[3671] =  13'b0000110100001; // 417 0.10173363238573074
storage[3672] =  13'b0000010110001; // 177 0.04331165552139282
storage[3673] =  13'b0000000011000; // 24 0.005916147492825985
storage[3674] = -13'b0000010111111; // -191 -0.046640921384096146
storage[3675] = -13'b0000001011110; // -94 -0.02299400232732296
storage[3676] =  13'b0000000000111; // 7 0.001805549836717546
storage[3677] = -13'b0000001110101; // -117 -0.02854362688958645
storage[3678] = -13'b0000011111100; // -252 -0.0616433210670948
storage[3679] =  13'b0000010001111; // 143 0.03496025502681732
storage[3680] = -13'b0000000101111; // -47 -0.011488568037748337
storage[3681] =  13'b0000010110001; // 177 0.04330841079354286
storage[3682] = -13'b0000000011100; // -28 -0.006919506471604109
storage[3683] = -13'b0000010101010; // -170 -0.04162066429853439
storage[3684] = -13'b0001001001001; // -585 -0.14282551407814026
storage[3685] = -13'b0000011000001; // -193 -0.04709810018539429
storage[3686] = -13'b0000000100110; // -38 -0.009378907270729542
storage[3687] = -13'b0000001111011; // -123 -0.029988018795847893
storage[3688] = -13'b0000000001001; // -9 -0.0021740002557635307
storage[3689] = -13'b0000001011111; // -95 -0.023132795467972755
storage[3690] = -13'b0000001110110; // -118 -0.02878670021891594
storage[3691] = -13'b0000001101011; // -107 -0.026118449866771698
storage[3692] =  13'b0000010011111; // 159 0.038878317922353745
storage[3693] =  13'b0000011111010; // 250 0.06105528399348259
storage[3694] =  13'b0000000111011; // 59 0.014282514341175556
storage[3695] = -13'b0000101101000; // -360 -0.08798031508922577
storage[3696] =  13'b0000010001011; // 139 0.0338367335498333
storage[3697] = -13'b0000010000110; // -134 -0.03276141732931137
storage[3698] =  13'b0000001011111; // 95 0.0232195183634758
storage[3699] =  13'b0000101000000; // 320 0.07820111513137817
storage[3700] = -13'b0000011110001; // -241 -0.05872909724712372
storage[3701] =  13'b0001001000000; // 576 0.14059039950370789
storage[3702] = -13'b0000100101010; // -298 -0.07275371253490448
storage[3703] =  13'b0000100100010; // 290 0.070711150765419
storage[3704] =  13'b0010010111111; // 1215 0.296749085187912
storage[3705] =  13'b0000110000011; // 387 0.09457747638225555
storage[3706] = -13'b0000001001111; // -79 -0.01935500279068947
storage[3707] = -13'b0000101111000; // -376 -0.09185129404067993
storage[3708] = -13'b0000000001000; // -8 -0.002070003654807806
storage[3709] =  13'b0000110100010; // 418 0.1021030992269516
storage[3710] =  13'b0001000010101; // 533 0.13018940389156342
storage[3711] =  13'b0000010111011; // 187 0.0456351712346077
storage[3712] = -13'b0000100101001; // -297 -0.07256459444761276
storage[3713] = -13'b0001001101000; // -616 -0.15044839680194855
storage[3714] =  13'b0000000100111; // 39 0.00952588114887476
storage[3715] = -13'b0000100111011; // -315 -0.07695110142230988
storage[3716] = -13'b0000111011100; // -476 -0.11627189069986343
storage[3717] =  13'b0000011111101; // 253 0.061775825917720795
storage[3718] = -13'b0000110111101; // -445 -0.10859330743551254
storage[3719] = -13'b0000011010100; // -212 -0.05164512246847153
storage[3720] =  13'b0000001111110; // 126 0.030725345015525818
storage[3721] =  13'b0000001000000; // 64 0.015597304329276085
storage[3722] = -13'b0000000101110; // -46 -0.011316077783703804
storage[3723] = -13'b0000001101010; // -106 -0.025870108976960182
storage[3724] =  13'b0000000110101; // 53 0.012849239632487297
storage[3725] =  13'b0000001100000; // 96 0.02353070303797722
storage[3726] = -13'b0001000101100; // -556 -0.135652557015419
storage[3727] = -13'b0000011001100; // -204 -0.04969006031751633
storage[3728] = -13'b0000111100110; // -486 -0.11858478933572769
storage[3729] = -13'b0001001101011; // -619 -0.15108726918697357
storage[3730] = -13'b0000011101111; // -239 -0.05845062807202339
storage[3731] = -13'b0000110000111; // -391 -0.09555098414421082
storage[3732] = -13'b0000011101101; // -237 -0.05779552832245827
storage[3733] = -13'b0000101001010; // -330 -0.08066194504499435
storage[3734] = -13'b0001010110111; // -695 -0.16958875954151154
storage[3735] = -13'b0000001011001; // -89 -0.021824663504958153
storage[3736] =  13'b0000011010000; // 208 0.05070647597312927
storage[3737] =  13'b0000011001101; // 205 0.050003983080387115
storage[3738] =  13'b0000010110101; // 181 0.04423262178897858
storage[3739] = -13'b0000001110001; // -113 -0.027529938146471977
storage[3740] = -13'b0000010111010; // -186 -0.04544871300458908
storage[3741] = -13'b0000001000001; // -65 -0.015769382938742638
storage[3742] =  13'b0000000001000; // 8 0.0020350904669612646
storage[3743] = -13'b0000011000011; // -195 -0.04768941551446915
storage[3744] = -13'b0000000001110; // -14 -0.0034314822405576706
storage[3745] = -13'b0000111011011; // -475 -0.11601495742797852
storage[3746] = -13'b0000010000110; // -134 -0.03278821334242821
storage[3747] =  13'b0000010000111; // 135 0.033030278980731964
storage[3748] = -13'b0000010101111; // -175 -0.04279058799147606
storage[3749] = -13'b0000101001100; // -332 -0.08105640858411789
storage[3750] = -13'b0000100101000; // -296 -0.07215369492769241
storage[3751] =  13'b0000110001001; // 393 0.09606669843196869
storage[3752] =  13'b0001001001111; // 591 0.14421528577804565
storage[3753] = -13'b0000000111010; // -58 -0.014163034968078136
storage[3754] = -13'b0000001001100; // -76 -0.018537301570177078
storage[3755] =  13'b0000100110111; // 311 0.0760296881198883
storage[3756] =  13'b0000001100011; // 99 0.02408606931567192
storage[3757] =  13'b0000001101010; // 106 0.025923142209649086
storage[3758] = -13'b0000011001110; // -206 -0.05031328275799751
storage[3759] = -13'b0000011100110; // -230 -0.05607268959283829
storage[3760] =  13'b0000011000001; // 193 0.04700084775686264
storage[3761] = -13'b0000101001101; // -333 -0.08136259764432907
storage[3762] = -13'b0000000110110; // -54 -0.013148502446711063
storage[3763] = -13'b0000101011011; // -347 -0.08481067419052124
storage[3764] =  13'b0000010001001; // 137 0.03334438428282738
storage[3765] =  13'b0000100011001; // 281 0.06863657385110855
storage[3766] = -13'b0001010111110; // -702 -0.17128148674964905
storage[3767] = -13'b0000010100111; // -167 -0.04083671420812607
storage[3768] = -13'b0000101100000; // -352 -0.08604110032320023
storage[3769] =  13'b0000011011010; // 218 0.05318927392363548
storage[3770] =  13'b0000110000110; // 390 0.0951419547200203
storage[3771] = -13'b0000010000111; // -135 -0.0329759307205677
storage[3772] =  13'b0000001010111; // 87 0.021249622106552124
storage[3773] =  13'b0000001110100; // 116 0.028430430218577385
storage[3774] = -13'b0000000000100; // -4 -0.0009284242987632751
storage[3775] =  13'b0000100010111; // 279 0.06822519749403
storage[3776] = -13'b0000000011010; // -26 -0.0062321326695382595
storage[3777] = -13'b0000010011011; // -155 -0.03786187991499901
storage[3778] =  13'b0000011011000; // 216 0.052612874656915665
storage[3779] =  13'b0000100010101; // 277 0.06763049215078354
storage[3780] =  13'b0000100111110; // 318 0.0777401551604271
storage[3781] =  13'b0000010010011; // 147 0.035941243171691895
storage[3782] =  13'b0000011000000; // 192 0.04685487970709801
storage[3783] =  13'b0000000011011; // 27 0.006526122335344553
storage[3784] = -13'b0000000101100; // -44 -0.010779895819723606
storage[3785] = -13'b0000100001111; // -271 -0.06607107073068619
storage[3786] = -13'b0000100101011; // -299 -0.07303030788898468
storage[3787] = -13'b0000010001101; // -141 -0.0344119630753994
storage[3788] =  13'b0000101101111; // 367 0.08960164338350296
storage[3789] =  13'b0000110110111; // 439 0.10711154341697693
storage[3790] = -13'b0001000000101; // -517 -0.12619082629680634
storage[3791] = -13'b0000110001111; // -399 -0.09748035669326782
storage[3792] =  13'b0000010100000; // 160 0.03906732797622681
storage[3793] = -13'b0000000011100; // -28 -0.006728159263730049
storage[3794] =  13'b0000010011100; // 156 0.038011111319065094
storage[3795] = -13'b0000011000010; // -194 -0.04729306325316429
storage[3796] =  13'b0000001000111; // 71 0.01738079823553562
storage[3797] =  13'b0000111110011; // 499 0.12180919945240021
storage[3798] =  13'b0000011000111; // 199 0.048632510006427765
storage[3799] = -13'b0000000101000; // -40 -0.009672936983406544
storage[3800] =  13'b0000110110011; // 435 0.10617314279079437
storage[3801] =  13'b0000001100001; // 97 0.023591144010424614
storage[3802] = -13'b0000101001100; // -332 -0.08095769584178925
storage[3803] =  13'b0001000100110; // 550 0.13433076441287994
storage[3804] =  13'b0000011100000; // 224 0.05456947535276413
storage[3805] =  13'b0000000110111; // 55 0.013549469411373138
storage[3806] =  13'b0000001011101; // 93 0.022695938125252724
storage[3807] =  13'b0000001010100; // 84 0.02048259787261486
storage[3808] = -13'b0000001100011; // -99 -0.02411300130188465
storage[3809] = -13'b0000101110000; // -368 -0.0899280235171318
storage[3810] =  13'b0000001001100; // 76 0.01866198144853115
storage[3811] =  13'b0000000001111; // 15 0.003561410354450345
storage[3812] =  13'b0000000010100; // 20 0.0049988445825874805
storage[3813] = -13'b0000001101001; // -105 -0.02560386061668396
storage[3814] = -13'b0000100011001; // -281 -0.06850948184728622
storage[3815] = -13'b0001111000100; // -964 -0.23540857434272766
storage[3816] = -13'b0000001111100; // -124 -0.030305197462439537
storage[3817] = -13'b0001100100011; // -803 -0.19610366225242615
storage[3818] = -13'b0000110110000; // -432 -0.10537069290876389
storage[3819] = -13'b0000100110011; // -307 -0.07503733783960342
storage[3820] = -13'b0001001011011; // -603 -0.14713986217975616
storage[3821] = -13'b0000101100010; // -354 -0.08654610067605972
storage[3822] =  13'b0000001010000; // 80 0.01964898407459259
storage[3823] = -13'b0001010011001; // -665 -0.16236019134521484
storage[3824] =  13'b0000001000101; // 69 0.016884319484233856
storage[3825] =  13'b0000100010011; // 275 0.06720443814992905
storage[3826] =  13'b0000000001001; // 9 0.00222381460480392
storage[3827] =  13'b0000010010110; // 150 0.03654203191399574
storage[3828] = -13'b0001001001011; // -587 -0.14333654940128326
storage[3829] = -13'b0000010011100; // -156 -0.03806636109948158
storage[3830] =  13'b0000100110010; // 306 0.07473262399435043
storage[3831] =  13'b0000100111110; // 318 0.07774651795625687
storage[3832] = -13'b0000010101110; // -174 -0.042410969734191895
storage[3833] =  13'b0000000110111; // 55 0.013369474560022354
storage[3834] =  13'b0000001000000; // 64 0.015690797939896584
storage[3835] =  13'b0000100110001; // 305 0.07454876601696014
storage[3836] =  13'b0000011100001; // 225 0.05487519130110741
storage[3837] = -13'b0000101101010; // -362 -0.08846651017665863
storage[3838] =  13'b0000101100101; // 357 0.08723780512809753
storage[3839] =  13'b0001000001101; // 525 0.12817290425300598
storage[3840] =  13'b0000000110101; // 53 0.013055999763309956
storage[3841] =  13'b0000100001011; // 267 0.06522540748119354
storage[3842] =  13'b0000010101001; // 169 0.0412178672850132
storage[3843] =  13'b0000100110110; // 310 0.07577618211507797
storage[3844] = -13'b0000110011001; // -409 -0.09991457313299179
storage[3845] =  13'b0000011001111; // 207 0.05055120587348938
storage[3846] =  13'b0000011001111; // 207 0.05059589445590973
storage[3847] = -13'b0000100010011; // -275 -0.06723611801862717
storage[3848] =  13'b0000000110010; // 50 0.012256978079676628
storage[3849] =  13'b0000001100011; // 99 0.024251513183116913
storage[3850] =  13'b0000001001110; // 78 0.019030818715691566
storage[3851] = -13'b0000001110000; // -112 -0.027433933690190315
storage[3852] =  13'b0000101101011; // 363 0.08855780959129333
storage[3853] = -13'b0000110010001; // -401 -0.09781957417726517
storage[3854] =  13'b0000011100101; // 229 0.05580532178282738
storage[3855] =  13'b0001000100110; // 550 0.13432075083255768
storage[3856] = -13'b0000010101001; // -169 -0.04118938744068146
storage[3857] =  13'b0000000100111; // 39 0.009557707235217094
storage[3858] =  13'b0000011111110; // 254 0.06206193566322327
storage[3859] =  13'b0000000011100; // 28 0.0067672329023480415
storage[3860] =  13'b0000010111001; // 185 0.045086268335580826
storage[3861] =  13'b0001001010100; // 596 0.1455061137676239
storage[3862] =  13'b0000000001001; // 9 0.0023042866960167885
storage[3863] = -13'b0000001000011; // -67 -0.016441121697425842
storage[3864] = -13'b0000001100100; // -100 -0.024302169680595398
storage[3865] = -13'b0000001110000; // -112 -0.02743816375732422
storage[3866] = -13'b0000111110100; // -500 -0.12201960384845734
storage[3867] = -13'b0000010010111; // -151 -0.03683847188949585
storage[3868] =  13'b0000011100110; // 230 0.05619170516729355
storage[3869] =  13'b0000100000010; // 258 0.06310760229825974
storage[3870] =  13'b0000100100100; // 292 0.07127483189105988
storage[3871] = -13'b0000001010111; // -87 -0.02131018415093422
storage[3872] = -13'b0000010010110; // -150 -0.03657519444823265
storage[3873] = -13'b0000101100111; // -359 -0.08754298835992813
storage[3874] = -13'b0001000000110; // -518 -0.12636218965053558
storage[3875] = -13'b0001111001111; // -975 -0.23801082372665405
storage[3876] = -13'b0000000011100; // -28 -0.006916950456798077
storage[3877] = -13'b0001111111110; // -1022 -0.24961689114570618
storage[3878] = -13'b0000101111011; // -379 -0.09241727739572525
storage[3879] =  13'b0000011011011; // 219 0.05343668535351753
storage[3880] = -13'b0000001110101; // -117 -0.02859220653772354
storage[3881] =  13'b0000000110101; // 53 0.012896944768726826
storage[3882] = -13'b0000000100000; // -32 -0.007794314529746771
storage[3883] =  13'b0000001011000; // 88 0.021423276513814926
storage[3884] =  13'b0000001111010; // 122 0.029906723648309708
storage[3885] = -13'b0000011010100; // -212 -0.051776304841041565
storage[3886] = -13'b0000011011011; // -219 -0.053526706993579865
storage[3887] = -13'b0000000001010; // -10 -0.0024012718349695206
storage[3888] =  13'b0000110000101; // 389 0.0948529839515686
storage[3889] = -13'b0000100001100; // -268 -0.06544409692287445
storage[3890] = -13'b0000100011110; // -286 -0.06985670328140259
storage[3891] = -13'b0000100011000; // -280 -0.06837178766727448
storage[3892] =  13'b0000110001010; // 394 0.0962720587849617
storage[3893] =  13'b0000001111100; // 124 0.030330467969179153
storage[3894] =  13'b0000011101110; // 238 0.05815032869577408
storage[3895] = -13'b0000000000010; // -2 -0.00044364179484546185
storage[3896] = -13'b0000010011000; // -152 -0.03719128668308258
storage[3897] = -13'b0000001000001; // -65 -0.015883907675743103
storage[3898] = -13'b0000000110101; // -53 -0.013013939373195171
storage[3899] = -13'b0000001110011; // -115 -0.027974506840109825
storage[3900] =  13'b0000000111111; // 63 0.01538895070552826
storage[3901] = -13'b0000110111001; // -441 -0.10755714774131775
storage[3902] = -13'b0000011010101; // -213 -0.05192447081208229
storage[3903] =  13'b0000011010000; // 208 0.05075763911008835
storage[3904] =  13'b0000001101111; // 111 0.02715563029050827
storage[3905] =  13'b0000101000100; // 324 0.07900784909725189
storage[3906] =  13'b0000100100111; // 295 0.0719560831785202
storage[3907] =  13'b0000110110010; // 434 0.10600442439317703
storage[3908] =  13'b0000101010001; // 337 0.08219877630472183
storage[3909] =  13'b0000110100001; // 417 0.10191088169813156
storage[3910] =  13'b0000101100000; // 352 0.0858229249715805
storage[3911] =  13'b0000101101000; // 360 0.08791696280241013
storage[3912] = -13'b0000100010100; // -276 -0.0673704594373703
storage[3913] = -13'b0000100010100; // -276 -0.06730122864246368
storage[3914] =  13'b0000100001110; // 270 0.06593132019042969
storage[3915] = -13'b0000001011001; // -89 -0.021614843979477882
storage[3916] = -13'b0001011010100; // -724 -0.176763117313385
storage[3917] = -13'b0000000011001; // -25 -0.006201264448463917
storage[3918] =  13'b0000001000010; // 66 0.01618589647114277
storage[3919] = -13'b0000001001100; // -76 -0.018630212172865868
storage[3920] = -13'b0000000100110; // -38 -0.009304944425821304
storage[3921] = -13'b0001000001111; // -527 -0.12875787913799286
storage[3922] = -13'b0000001100010; // -98 -0.023885389789938927
storage[3923] = -13'b0000110001101; // -397 -0.09702790528535843
storage[3924] = -13'b0001000011000; // -536 -0.1308794915676117
storage[3925] = -13'b0000111010100; // -468 -0.1142827644944191
storage[3926] =  13'b0000001100110; // 102 0.024977752938866615
storage[3927] =  13'b0000101101111; // 367 0.08964324742555618
storage[3928] = -13'b0001101001001; // -841 -0.20523594319820404
storage[3929] =  13'b0000010111100; // 188 0.0458604097366333
storage[3930] =  13'b0000011010000; // 208 0.05083424225449562
storage[3931] = -13'b0000111110101; // -501 -0.12230665981769562
storage[3932] =  13'b0000000001000; // 8 0.0019585243426263332
storage[3933] =  13'b0000011010101; // 213 0.05205807834863663
storage[3934] =  13'b0001000100100; // 548 0.13372613489627838
storage[3935] =  13'b0000011001101; // 205 0.04996674135327339
storage[3936] =  13'b0000001000000; // 64 0.015507019124925137
storage[3937] = -13'b0000000110011; // -51 -0.012448441237211227
storage[3938] =  13'b0000001011100; // 92 0.022347381338477135
storage[3939] =  13'b0000001100001; // 97 0.02365581877529621
storage[3940] = -13'b0000000000000; // 0 -0.0001067309349309653
storage[3941] = -13'b0000000101101; // -45 -0.010887826792895794
storage[3942] =  13'b0000001101111; // 111 0.027084028348326683
storage[3943] =  13'b0000000011111; // 31 0.0074781919829547405
storage[3944] = -13'b0000100110101; // -309 -0.07534634321928024
storage[3945] = -13'b0001001000011; // -579 -0.14123719930648804
storage[3946] =  13'b0000010100110; // 166 0.040597155690193176
storage[3947] = -13'b0000010001011; // -139 -0.03387495130300522
storage[3948] = -13'b0000101010011; // -339 -0.08264379948377609
storage[3949] =  13'b0000010111110; // 190 0.04645884782075882
storage[3950] = -13'b0000010111111; // -191 -0.046596772968769073
storage[3951] =  13'b0000001011011; // 91 0.02221526764333248
storage[3952] = -13'b0000000001101; // -13 -0.003162339562550187
storage[3953] =  13'b0000001111111; // 127 0.03110477514564991
storage[3954] =  13'b0000100001101; // 269 0.06561906635761261
storage[3955] =  13'b0000000110000; // 48 0.011699614115059376
storage[3956] =  13'b0000001110101; // 117 0.02859725058078766
storage[3957] =  13'b0000011101101; // 237 0.05785737931728363
storage[3958] =  13'b0000000010011; // 19 0.004555744584649801
storage[3959] =  13'b0000100110101; // 309 0.07555745542049408
storage[3960] =  13'b0000100000001; // 257 0.06264913082122803
storage[3961] =  13'b0000110000110; // 390 0.095257967710495
storage[3962] =  13'b0000001001011; // 75 0.018211379647254944
storage[3963] =  13'b0000011111100; // 252 0.061502452939748764
storage[3964] =  13'b0000001011000; // 88 0.021566519513726234
storage[3965] = -13'b0000000001000; // -8 -0.0019730492495000362
storage[3966] = -13'b0000000001110; // -14 -0.0034825389739125967
storage[3967] =  13'b0000000010110; // 22 0.005345530807971954
storage[3968] =  13'b0000011101110; // 238 0.05820292979478836
storage[3969] =  13'b0000100011011; // 283 0.06916237622499466
storage[3970] = -13'b0000110001100; // -396 -0.09672722220420837
storage[3971] = -13'b0000010111011; // -187 -0.04575423523783684
storage[3972] =  13'b0000001100111; // 103 0.02519724890589714
storage[3973] = -13'b0000101100000; // -352 -0.08593863993883133
storage[3974] = -13'b0000001000111; // -71 -0.01735992543399334
storage[3975] =  13'b0000010010111; // 151 0.03676123917102814
storage[3976] =  13'b0000110011111; // 415 0.10135629773139954
storage[3977] =  13'b0000101010110; // 342 0.08345480263233185
storage[3978] =  13'b0000101111000; // 376 0.09187203645706177
storage[3979] =  13'b0000010100101; // 165 0.04032120481133461
storage[3980] =  13'b0000000010010; // 18 0.004471180960536003
storage[3981] =  13'b0000000001101; // 13 0.003282850841060281
storage[3982] =  13'b0000100001100; // 268 0.0653373971581459
storage[3983] =  13'b0000000100111; // 39 0.009486613795161247
storage[3984] = -13'b0000100000000; // -256 -0.06247150897979736
storage[3985] = -13'b0000000101101; // -45 -0.010873612947762012
storage[3986] =  13'b0000001111000; // 120 0.029294423758983612
storage[3987] =  13'b0000011101000; // 232 0.05652236565947533
storage[3988] = -13'b0000010101011; // -171 -0.04165124520659447
storage[3989] =  13'b0000011011100; // 220 0.05366719514131546
storage[3990] = -13'b0000011110010; // -242 -0.059159304946660995
storage[3991] =  13'b0000000110100; // 52 0.012585317716002464
storage[3992] =  13'b0000100001011; // 267 0.06520187854766846
storage[3993] = -13'b0000000101011; // -43 -0.010569017380475998
storage[3994] =  13'b0000011001101; // 205 0.05012763291597366
storage[3995] =  13'b0000000110011; // 51 0.012364529073238373
storage[3996] =  13'b0000010100001; // 161 0.03930521383881569
storage[3997] =  13'b0000001100000; // 96 0.023349102586507797
storage[3998] =  13'b0000000010000; // 16 0.003810859750956297
storage[3999] = -13'b0000000010101; // -21 -0.00509868748486042
storage[4000] =  13'b0000000010100; // 20 0.004843195900321007
storage[4001] =  13'b0000001001001; // 73 0.01793205551803112
storage[4002] =  13'b0000000110110; // 54 0.013080721721053123
storage[4003] =  13'b0000001110011; // 115 0.027964157983660698
storage[4004] = -13'b0000001101010; // -106 -0.02596011944115162
storage[4005] = -13'b0000010000100; // -132 -0.03224428370594978
storage[4006] =  13'b0000000111000; // 56 0.013654245994985104
storage[4007] =  13'b0000000111000; // 56 0.013653668574988842
storage[4008] = -13'b0000011001101; // -205 -0.05013403668999672
storage[4009] = -13'b0000011001110; // -206 -0.0503111332654953
storage[4010] =  13'b0000100010100; // 276 0.06729058921337128
storage[4011] =  13'b0000001010010; // 82 0.020088056102395058
storage[4012] = -13'b0000011000101; // -197 -0.048029229044914246
storage[4013] =  13'b0000100110011; // 307 0.07505927979946136
storage[4014] =  13'b0000100101111; // 303 0.0739300474524498
storage[4015] = -13'b0000110001000; // -392 -0.0957338884472847
storage[4016] = -13'b0000001001011; // -75 -0.01825217343866825
storage[4017] =  13'b0000010111011; // 187 0.04570163041353226
storage[4018] = -13'b0000010000010; // -130 -0.03170393407344818
storage[4019] = -13'b0000000000001; // -1 -0.0002897191734518856
storage[4020] = -13'b0000011101000; // -232 -0.05652054771780968
storage[4021] = -13'b0000100101111; // -303 -0.07393713295459747
storage[4022] =  13'b0000000011000; // 24 0.005873213522136211
storage[4023] = -13'b0000001001111; // -79 -0.019178763031959534
storage[4024] = -13'b0000001110000; // -112 -0.027453593909740448
storage[4025] =  13'b0001100111101; // 829 0.20245492458343506
storage[4026] =  13'b0000001001011; // 75 0.018352866172790527
storage[4027] = -13'b0000101110001; // -369 -0.08998818695545197
storage[4028] = -13'b0001000100110; // -550 -0.13423112034797668
storage[4029] =  13'b0000000011011; // 27 0.006627578753978014
storage[4030] = -13'b0000001011100; // -92 -0.022579442709684372
storage[4031] = -13'b0001001101110; // -622 -0.15184657275676727
storage[4032] = -13'b0000111110001; // -497 -0.12137538194656372
storage[4033] =  13'b0000000110011; // 51 0.012517409399151802
storage[4034] = -13'b0001001011000; // -600 -0.14640095829963684
storage[4035] = -13'b0000110101000; // -424 -0.10344894230365753
storage[4036] =  13'b0000100001101; // 269 0.0656515583395958
storage[4037] =  13'b0000001011001; // 89 0.0217672660946846
storage[4038] =  13'b0000010000011; // 131 0.0320102721452713
storage[4039] =  13'b0000100110001; // 305 0.07441068440675735
storage[4040] = -13'b0000011010100; // -212 -0.05174606293439865
storage[4041] =  13'b0000010100111; // 167 0.040725573897361755
storage[4042] =  13'b0000110111010; // 442 0.10796989500522614
storage[4043] =  13'b0000010000101; // 133 0.03249521180987358
storage[4044] =  13'b0000011110010; // 242 0.059189822524785995
storage[4045] =  13'b0000001101111; // 111 0.026994772255420685
storage[4046] = -13'b0000100000001; // -257 -0.06281010061502457
storage[4047] =  13'b0000110100010; // 418 0.10201582312583923
storage[4048] =  13'b0000101000000; // 320 0.07811354100704193
storage[4049] = -13'b0000000101010; // -42 -0.010247698985040188
storage[4050] =  13'b0001001100100; // 612 0.14948734641075134
storage[4051] =  13'b0000000111110; // 62 0.01517743244767189
storage[4052] = -13'b0000001101010; // -106 -0.0258793905377388
storage[4053] = -13'b0000101010000; // -336 -0.08210182934999466
storage[4054] =  13'b0000110000001; // 385 0.09393687546253204
storage[4055] =  13'b0000001010111; // 87 0.021124260500073433
storage[4056] =  13'b0000001011000; // 88 0.021388763561844826
storage[4057] = -13'b0000000110110; // -54 -0.013080505654215813
storage[4058] =  13'b0000011011000; // 216 0.05263160541653633
storage[4059] = -13'b0000001100001; // -97 -0.02358049899339676
storage[4060] =  13'b0000011001101; // 205 0.050102755427360535
storage[4061] =  13'b0000001101110; // 110 0.026973458006978035
storage[4062] = -13'b0000001100001; // -97 -0.0237205158919096
storage[4063] = -13'b0000000011001; // -25 -0.006154290866106749
storage[4064] =  13'b0000111110111; // 503 0.12288130074739456
storage[4065] =  13'b0000101110010; // 370 0.09022404253482819
storage[4066] =  13'b0000100100010; // 290 0.07072649896144867
storage[4067] =  13'b0001001001110; // 590 0.14397038519382477
storage[4068] =  13'b0000011000000; // 192 0.04688943922519684
storage[4069] = -13'b0000101110010; // -370 -0.09039246290922165
storage[4070] = -13'b0001001011011; // -603 -0.1472810059785843
storage[4071] = -13'b0000100110011; // -307 -0.07498753070831299
storage[4072] =  13'b0000100101100; // 300 0.0732017531991005
storage[4073] = -13'b0000001110001; // -113 -0.027605580165982246
storage[4074] = -13'b0000000001111; // -15 -0.0035454921890050173
storage[4075] =  13'b0000001000101; // 69 0.01677563786506653
storage[4076] = -13'b0000001110110; // -118 -0.028742708265781403
storage[4077] =  13'b0000010000000; // 128 0.031303051859140396
storage[4078] = -13'b0001011111101; // -765 -0.18667858839035034
storage[4079] = -13'b0000111001110; // -462 -0.11267708241939545
storage[4080] = -13'b0001101001001; // -841 -0.20526383817195892
storage[4081] = -13'b0000000000110; // -6 -0.0015382893616333604
storage[4082] = -13'b0000001110010; // -114 -0.027847876772284508
storage[4083] = -13'b0000001110010; // -114 -0.027759015560150146
storage[4084] = -13'b0000010001011; // -139 -0.034055449068546295
storage[4085] =  13'b0000011100111; // 231 0.05631197616457939
storage[4086] =  13'b0000010100000; // 160 0.03910183906555176
storage[4087] =  13'b0000110001101; // 397 0.09699279069900513
storage[4088] =  13'b0001001000110; // 582 0.14212144911289215
storage[4089] = -13'b0000000001001; // -9 -0.0022003690246492624
storage[4090] =  13'b0000101011101; // 349 0.08527883887290955
storage[4091] =  13'b0000101000011; // 323 0.07877235114574432
storage[4092] =  13'b0000100001100; // 268 0.06547260284423828
storage[4093] = -13'b0000000100001; // -33 -0.008111714385449886
storage[4094] =  13'b0000110101010; // 426 0.10408143699169159
storage[4095] = -13'b0000010111110; // -190 -0.04635613411664963
storage[4096] = -13'b0000010011101; // -157 -0.0382971428334713
storage[4097] = -13'b0000001010111; // -87 -0.0213572196662426
storage[4098] =  13'b0000011100111; // 231 0.056357771158218384
storage[4099] = -13'b0000100110110; // -310 -0.07565666735172272
storage[4100] =  13'b0000000010111; // 23 0.005684655159711838
storage[4101] = -13'b0000010111011; // -187 -0.04566708952188492
storage[4102] =  13'b0000001100000; // 96 0.023459475487470627
storage[4103] =  13'b0000001100001; // 97 0.02371450699865818
storage[4104] = -13'b0000011010011; // -211 -0.05140788480639458
storage[4105] =  13'b0000010001000; // 136 0.033208854496479034
storage[4106] =  13'b0000010000111; // 135 0.03284215182065964
storage[4107] = -13'b0001000001000; // -520 -0.12685811519622803
storage[4108] =  13'b0000100000101; // 261 0.0637938603758812
storage[4109] =  13'b0000011101100; // 236 0.05756840109825134
storage[4110] = -13'b0000000101010; // -42 -0.010149587877094746
storage[4111] =  13'b0000010010000; // 144 0.03514830023050308
storage[4112] =  13'b0000101000100; // 324 0.07912459969520569
storage[4113] =  13'b0000010110101; // 181 0.0442175418138504
storage[4114] =  13'b0000000100111; // 39 0.00959260668605566
storage[4115] = -13'b0000011100111; // -231 -0.05643746629357338
storage[4116] = -13'b0000110011000; // -408 -0.09972374141216278
storage[4117] =  13'b0000001111110; // 126 0.03080267459154129
storage[4118] =  13'b0000000010101; // 21 0.005109262187033892
storage[4119] = -13'b0000001100011; // -99 -0.024219918996095657
storage[4120] =  13'b0000110100000; // 416 0.10144339501857758
storage[4121] =  13'b0000010011110; // 158 0.038612958043813705
storage[4122] =  13'b0000100110100; // 308 0.07509363442659378
storage[4123] = -13'b0000011111001; // -249 -0.06088534742593765
storage[4124] =  13'b0000001101101; // 109 0.026629682630300522
storage[4125] = -13'b0001010010010; // -658 -0.1606593132019043
storage[4126] = -13'b0000001000001; // -65 -0.015986748039722443
storage[4127] =  13'b0000010101100; // 172 0.04209836199879646
storage[4128] = -13'b0000110011111; // -415 -0.10120018571615219
storage[4129] =  13'b0000011010010; // 210 0.051165081560611725
storage[4130] =  13'b0000001101111; // 111 0.02708963118493557
storage[4131] =  13'b0000101101110; // 366 0.0893239974975586
storage[4132] = -13'b0000010011001; // -153 -0.037279654294252396
storage[4133] = -13'b0000000001101; // -13 -0.00326199596747756
storage[4134] =  13'b0000101011111; // 351 0.08557182550430298
storage[4135] = -13'b0000000101010; // -42 -0.010180734097957611
storage[4136] = -13'b0000000111010; // -58 -0.01428096741437912
storage[4137] = -13'b0000001110110; // -118 -0.02880486473441124
storage[4138] = -13'b0000010001001; // -137 -0.0335422158241272
storage[4139] = -13'b0000101100001; // -353 -0.08607754111289978
storage[4140] = -13'b0000010101010; // -170 -0.04162446781992912
storage[4141] = -13'b0000011111100; // -252 -0.06155781447887421
storage[4142] =  13'b0000011001110; // 206 0.05028662830591202
storage[4143] =  13'b0000010100010; // 162 0.039433106780052185
storage[4144] = -13'b0000000001100; // -12 -0.002951906993985176
storage[4145] = -13'b0001110011101; // -925 -0.22574114799499512
storage[4146] = -13'b0000010100101; // -165 -0.04040224105119705
storage[4147] =  13'b0000101111111; // 383 0.09361007809638977
storage[4148] =  13'b0000010010101; // 149 0.03632641211152077
storage[4149] =  13'b0000101001010; // 330 0.08063673228025436
storage[4150] = -13'b0000001111100; // -124 -0.030290769413113594
storage[4151] =  13'b0001010110001; // 689 0.16833117604255676
storage[4152] = -13'b0000101010000; // -336 -0.08206922560930252
storage[4153] =  13'b0000100110110; // 310 0.07571963220834732
storage[4154] =  13'b0000100111000; // 312 0.07616935670375824
storage[4155] = -13'b0000110010101; // -405 -0.09880868345499039
storage[4156] =  13'b0000000101100; // 44 0.010831876657903194
storage[4157] = -13'b0000100111010; // -314 -0.07673081755638123
storage[4158] = -13'b0001010000111; // -647 -0.15805339813232422
storage[4159] = -13'b0000110010110; // -406 -0.09923531115055084
storage[4160] = -13'b0000110100100; // -420 -0.102579265832901
storage[4161] = -13'b0000011010001; // -209 -0.051120661199092865
storage[4162] = -13'b0000110101101; // -429 -0.1048300713300705
storage[4163] = -13'b0000001010111; // -87 -0.02121444046497345
storage[4164] =  13'b0000000100011; // 35 0.008586296811699867
storage[4165] =  13'b0000011100111; // 231 0.05648915842175484
storage[4166] =  13'b0000001101000; // 104 0.025486774742603302
storage[4167] =  13'b0000100110001; // 305 0.07439998537302017
storage[4168] =  13'b0000010100011; // 163 0.039778657257556915
storage[4169] =  13'b0000000000110; // 6 0.0014879894442856312
storage[4170] = -13'b0001110100001; // -929 -0.22685228288173676
storage[4171] =  13'b0000100011011; // 283 0.06899083405733109
storage[4172] = -13'b0001000100010; // -546 -0.13340803980827332
storage[4173] = -13'b0000101110111; // -375 -0.09151682257652283
storage[4174] =  13'b0000100010101; // 277 0.06761519610881805
storage[4175] =  13'b0000000011100; // 28 0.006771288812160492
storage[4176] =  13'b0000000010100; // 20 0.004845269490033388
storage[4177] =  13'b0000111101010; // 490 0.11966709792613983
storage[4178] =  13'b0000000101000; // 40 0.009770127013325691
storage[4179] = -13'b0001010110101; // -693 -0.1691237986087799
storage[4180] =  13'b0000011000000; // 192 0.04684450104832649
storage[4181] =  13'b0000110100001; // 417 0.10176239162683487
storage[4182] =  13'b0000111001010; // 458 0.1118173748254776
storage[4183] =  13'b0000010110000; // 176 0.04306874796748161
storage[4184] =  13'b0000110011001; // 409 0.09993904829025269
storage[4185] =  13'b0000111100110; // 486 0.11869411170482635
storage[4186] =  13'b0000101011111; // 351 0.08575380593538284
storage[4187] =  13'b0000011111011; // 251 0.06129959970712662
storage[4188] = -13'b0000010010011; // -147 -0.03595948964357376
storage[4189] =  13'b0000110001001; // 393 0.09584149718284607
storage[4190] = -13'b0000111010101; // -469 -0.11451365053653717
storage[4191] =  13'b0001011011101; // 733 0.17888323962688446
storage[4192] = -13'b0000000010110; // -22 -0.0054154968820512295
storage[4193] = -13'b0001000101101; // -557 -0.13598312437534332
storage[4194] =  13'b0001101010000; // 848 0.20697082579135895
storage[4195] =  13'b0000011011010; // 218 0.05329286679625511
storage[4196] =  13'b0000001010001; // 81 0.01968081295490265
storage[4197] = -13'b0001001100011; // -611 -0.14919635653495789
storage[4198] =  13'b0000011000101; // 197 0.0480080246925354
storage[4199] = -13'b0000011000001; // -193 -0.047099366784095764
storage[4200] = -13'b0001110011001; // -921 -0.22496378421783447
storage[4201] =  13'b0000010001001; // 137 0.03350301459431648
storage[4202] = -13'b0000110001101; // -397 -0.09681317210197449
storage[4203] = -13'b0000011100011; // -227 -0.05552178993821144
storage[4204] =  13'b0000101100000; // 352 0.08604654669761658
storage[4205] =  13'b0000000001101; // 13 0.0031518612522631884
storage[4206] = -13'b0000100110110; // -310 -0.07579956948757172
storage[4207] =  13'b0000010011001; // 153 0.03744705766439438
storage[4208] = -13'b0010111011011; // -1499 -0.36602598428726196
storage[4209] = -13'b0000000110110; // -54 -0.013283479027450085
storage[4210] =  13'b0000101010011; // 339 0.08276648074388504
storage[4211] = -13'b0010000111100; // -1084 -0.2645968496799469
storage[4212] =  13'b0000110010111; // 407 0.09931116551160812
storage[4213] =  13'b0000010001011; // 139 0.03387649357318878
storage[4214] =  13'b0000010010011; // 147 0.03592405468225479
storage[4215] = -13'b0000001001001; // -73 -0.017802737653255463
storage[4216] = -13'b0000000000111; // -7 -0.0016932172002270818
storage[4217] = -13'b0000100001110; // -270 -0.06594580411911011
storage[4218] = -13'b0000000000001; // -1 -0.00021204260701779276
storage[4219] = -13'b0000001111001; // -121 -0.029624078422784805
storage[4220] =  13'b0000000101111; // 47 0.011398435570299625
storage[4221] = -13'b0000001001001; // -73 -0.017836356535553932
storage[4222] = -13'b0010000100011; // -1059 -0.25860798358917236
storage[4223] = -13'b0011010001110; // -1678 -0.40970534086227417
storage[4224] = -13'b0010000100011; // -1059 -0.25857749581336975
storage[4225] = -13'b0000101100101; // -357 -0.0871610939502716
storage[4226] = -13'b0000001101111; // -111 -0.027145126834511757
storage[4227] = -13'b0000101101011; // -363 -0.08855428546667099
storage[4228] =  13'b0000010111011; // 187 0.04561891779303551
storage[4229] =  13'b0000001000100; // 68 0.01669158786535263
storage[4230] =  13'b0000101000110; // 326 0.07963069528341293
storage[4231] =  13'b0000000011111; // 31 0.007652499713003635
storage[4232] = -13'b0000000110011; // -51 -0.012501206248998642
storage[4233] =  13'b0000010110010; // 178 0.04352673143148422
storage[4234] = -13'b0000000100000; // -32 -0.007879485376179218
storage[4235] =  13'b0000001101100; // 108 0.026383863762021065
storage[4236] =  13'b0000000110110; // 54 0.013189733028411865
storage[4237] =  13'b0000001000101; // 69 0.016757270321249962
storage[4238] =  13'b0000001001111; // 79 0.019167998805642128
storage[4239] = -13'b0000010000011; // -131 -0.03187970072031021
storage[4240] =  13'b0000001010110; // 86 0.021108917891979218
storage[4241] =  13'b0000001000010; // 66 0.016147350892424583
storage[4242] = -13'b0000001000101; // -69 -0.01696174032986164
storage[4243] =  13'b0000000111010; // 58 0.014276796951889992
storage[4244] =  13'b0000001111011; // 123 0.030015865340828896
storage[4245] =  13'b0000100000111; // 263 0.0642339438199997
storage[4246] =  13'b0000011101011; // 235 0.057385530322790146
storage[4247] =  13'b0000010011100; // 156 0.03811273351311684
storage[4248] = -13'b0000000110101; // -53 -0.012877973727881908
storage[4249] = -13'b0000100001000; // -264 -0.06447906792163849
storage[4250] =  13'b0000001101000; // 104 0.025459710508584976
storage[4251] = -13'b0000000000001; // -1 -0.00023639264691155404
storage[4252] =  13'b0000100110001; // 305 0.074351005256176
storage[4253] = -13'b0000000010111; // -23 -0.0055942232720553875
storage[4254] = -13'b0001100100100; // -804 -0.19621321558952332
storage[4255] = -13'b0000010010101; // -149 -0.036433134227991104
storage[4256] = -13'b0000100110110; // -310 -0.0756860226392746
storage[4257] = -13'b0000010101010; // -170 -0.04157666116952896
storage[4258] = -13'b0001000010001; // -529 -0.1291767656803131
storage[4259] = -13'b0000001011010; // -90 -0.021906791254878044
storage[4260] = -13'b0000000101110; // -46 -0.011275301687419415
storage[4261] =  13'b0000000111110; // 62 0.015135614201426506
storage[4262] =  13'b0000000011110; // 30 0.007352410349994898
storage[4263] = -13'b0010001011101; // -1117 -0.2727203667163849
storage[4264] =  13'b0000000101010; // 42 0.010280302725732327
storage[4265] = -13'b0000001110101; // -117 -0.028448564931750298
storage[4266] = -13'b0000100000101; // -261 -0.06364615261554718
storage[4267] = -13'b0001000101111; // -559 -0.13654205203056335
storage[4268] = -13'b0001011110101; // -757 -0.18473975360393524
storage[4269] =  13'b0000010110111; // 183 0.04471822455525398
storage[4270] = -13'b0000111000010; // -450 -0.10991901904344559
storage[4271] = -13'b0001011101111; // -751 -0.18324247002601624
storage[4272] = -13'b0001010000011; // -643 -0.15686753392219543
storage[4273] =  13'b0000101001010; // 330 0.08059521019458771
storage[4274] =  13'b0000110110000; // 432 0.10537704825401306
storage[4275] =  13'b0000110000100; // 388 0.0946163460612297
storage[4276] = -13'b0000000101100; // -44 -0.010713792406022549
storage[4277] = -13'b0000101000000; // -320 -0.07806069403886795
storage[4278] = -13'b0000000101001; // -41 -0.009963050484657288
storage[4279] = -13'b0000011000011; // -195 -0.047649215906858444
storage[4280] = -13'b0000011111010; // -250 -0.06113530322909355
storage[4281] = -13'b0000001001000; // -72 -0.017636427655816078
storage[4282] = -13'b0000100110000; // -304 -0.07427993416786194
storage[4283] =  13'b0000010111100; // 188 0.04585292190313339
storage[4284] =  13'b0000100001101; // 269 0.06563326716423035
storage[4285] = -13'b0000011011101; // -221 -0.053980376571416855
storage[4286] = -13'b0000011111100; // -252 -0.06146048381924629
storage[4287] = -13'b0000001110010; // -114 -0.027948962524533272
storage[4288] = -13'b0000011100100; // -228 -0.05572386458516121
storage[4289] =  13'b0000010110100; // 180 0.04384379833936691
storage[4290] =  13'b0000011000000; // 192 0.0467863455414772
storage[4291] =  13'b0000000001010; // 10 0.002370318863540888
storage[4292] =  13'b0000011101101; // 237 0.05775340273976326
storage[4293] =  13'b0000111011100; // 476 0.11615514010190964
storage[4294] =  13'b0000110001110; // 398 0.09716577082872391
storage[4295] = -13'b0000010110011; // -179 -0.043641168624162674
storage[4296] =  13'b0000000011100; // 28 0.006951770279556513
storage[4297] =  13'b0000111011110; // 478 0.11660480499267578
storage[4298] = -13'b0000010011001; // -153 -0.03737444058060646
storage[4299] =  13'b0000001011010; // 90 0.022056153044104576
storage[4300] =  13'b0001000011000; // 536 0.13096052408218384
storage[4301] =  13'b0000110011100; // 412 0.10047914832830429
storage[4302] = -13'b0000000000011; // -3 -0.0008157273405231535
storage[4303] = -13'b0000000001100; // -12 -0.0030452157370746136
storage[4304] =  13'b0000001110111; // 119 0.029121046885848045
storage[4305] =  13'b0000001111101; // 125 0.030523335561156273
storage[4306] = -13'b0000000000100; // -4 -0.0009433508384972811
storage[4307] = -13'b0000100000011; // -259 -0.06327849626541138
storage[4308] = -13'b0000101000111; // -327 -0.07982751727104187
storage[4309] = -13'b0000101000100; // -324 -0.07907746732234955
storage[4310] = -13'b0001000010110; // -534 -0.13047192990779877
storage[4311] = -13'b0000110101001; // -425 -0.10371514409780502
storage[4312] = -13'b0000011110011; // -243 -0.05929601937532425
storage[4313] = -13'b0000001011111; // -95 -0.023244867101311684
storage[4314] =  13'b0000101111000; // 376 0.09168127179145813
storage[4315] = -13'b0000011001100; // -204 -0.049711789935827255
storage[4316] = -13'b0001010011010; // -666 -0.16256925463676453
storage[4317] = -13'b0000011100111; // -231 -0.05642817169427872
storage[4318] = -13'b0000010001101; // -141 -0.03441851586103439
storage[4319] = -13'b0000110101010; // -426 -0.10405854135751724
storage[4320] = -13'b0000100001110; // -270 -0.06603357940912247
storage[4321] =  13'b0000011101010; // 234 0.05709782987833023
storage[4322] =  13'b0000001011011; // 91 0.022115077823400497
storage[4323] =  13'b0000011110010; // 242 0.059138793498277664
storage[4324] =  13'b0000000000010; // 2 0.0005540073616430163
storage[4325] = -13'b0000010001101; // -141 -0.0343211330473423
storage[4326] =  13'b0000100111110; // 318 0.07762744277715683
storage[4327] = -13'b0000001000001; // -65 -0.01579202152788639
storage[4328] = -13'b0000111000001; // -449 -0.10962271690368652
storage[4329] = -13'b0000011000100; // -196 -0.04789850860834122
storage[4330] =  13'b0000000000111; // 7 0.0016045988304540515
storage[4331] = -13'b0000100101000; // -296 -0.07235219329595566
storage[4332] = -13'b0000110101101; // -429 -0.10476861894130707
storage[4333] = -13'b0000011101101; // -237 -0.05793358385562897
storage[4334] = -13'b0000000011011; // -27 -0.006559509318321943
storage[4335] =  13'b0000000001111; // 15 0.0037018156144768
storage[4336] = -13'b0000011101110; // -238 -0.05818957835435867
storage[4337] = -13'b0000110011110; // -414 -0.1011543944478035
storage[4338] =  13'b0000001110101; // 117 0.02844688855111599
storage[4339] = -13'b0000010000100; // -132 -0.03219198063015938
storage[4340] = -13'b0000110011000; // -408 -0.09955006837844849
storage[4341] =  13'b0000001011010; // 90 0.021944602951407433
storage[4342] =  13'b0000100100000; // 288 0.07028844952583313
storage[4343] = -13'b0000000011111; // -31 -0.0076749371364712715
storage[4344] =  13'b0000110101010; // 426 0.10389461368322372
storage[4345] = -13'b0000000011111; // -31 -0.007643978111445904
storage[4346] = -13'b0000010010101; // -149 -0.036290302872657776
storage[4347] =  13'b0000000001000; // 8 0.0019992352463304996
storage[4348] = -13'b0000111101000; // -488 -0.11906951665878296
storage[4349] = -13'b0000011001011; // -203 -0.04944271221756935
storage[4350] = -13'b0000001111111; // -127 -0.031083162873983383
storage[4351] =  13'b0000011001011; // 203 0.049516547471284866
storage[4352] =  13'b0000011001011; // 203 0.04960716515779495
storage[4353] = -13'b0000100010011; // -275 -0.06709915399551392
storage[4354] = -13'b0000110011010; // -410 -0.10018337517976761
storage[4355] = -13'b0001101000000; // -832 -0.20321105420589447
storage[4356] = -13'b0001111110101; // -1013 -0.24736197292804718
storage[4357] =  13'b0000100010110; // 278 0.06779118627309799
storage[4358] = -13'b0000011111001; // -249 -0.06069951131939888
storage[4359] = -13'b0000101111001; // -377 -0.09215178340673447
storage[4360] =  13'b0000010000101; // 133 0.032578546553850174
storage[4361] =  13'b0000110000000; // 384 0.09365922212600708
storage[4362] =  13'b0000011110100; // 244 0.059492066502571106
storage[4363] =  13'b0000001100110; // 102 0.025021227076649666
storage[4364] =  13'b0000101010101; // 341 0.08320973068475723
storage[4365] =  13'b0000111001010; // 458 0.11172228306531906
storage[4366] =  13'b0000001010010; // 82 0.020111121237277985
storage[4367] =  13'b0000010111110; // 190 0.04650555178523064
storage[4368] =  13'b0000100010111; // 279 0.06814667582511902
storage[4369] =  13'b0000001001010; // 74 0.018132030963897705
storage[4370] =  13'b0001001000111; // 583 0.14224161207675934
storage[4371] =  13'b0000110000101; // 389 0.09492573887109756
storage[4372] =  13'b0000110011110; // 414 0.1011618971824646
storage[4373] =  13'b0000100010111; // 279 0.06820104271173477
storage[4374] = -13'b0000001100101; // -101 -0.024594267830252647
storage[4375] = -13'b0001000011010; // -538 -0.1312931627035141
storage[4376] = -13'b0000000110001; // -49 -0.012038064189255238
storage[4377] =  13'b0000000000011; // 3 0.0006216379697434604
storage[4378] = -13'b0000001100110; // -102 -0.02488187700510025
storage[4379] = -13'b0001000011100; // -540 -0.13188324868679047
storage[4380] =  13'b0000000011111; // 31 0.007677918765693903
storage[4381] = -13'b0000111000110; // -454 -0.11090906709432602
storage[4382] = -13'b0001000110001; // -561 -0.13699860870838165
storage[4383] = -13'b0000011111101; // -253 -0.06182783842086792
storage[4384] =  13'b0001001000011; // 579 0.1414109766483307
storage[4385] =  13'b0000001001011; // 75 0.01820238120853901
storage[4386] =  13'b0000000101110; // 46 0.011206446215510368
storage[4387] =  13'b0001000101111; // 559 0.13644765317440033
storage[4388] =  13'b0000100001110; // 270 0.06589225679636002
storage[4389] =  13'b0000010011011; // 155 0.037955768406391144
storage[4390] = -13'b0000010001101; // -141 -0.03446182236075401
storage[4391] = -13'b0000011100111; // -231 -0.05636383220553398
storage[4392] = -13'b0000110010010; // -402 -0.09816227108240128
storage[4393] = -13'b0000001100011; // -99 -0.02414979785680771
storage[4394] =  13'b0000001011001; // 89 0.021611331030726433
storage[4395] =  13'b0000000000000; // 0 3.71778583030391e-06
storage[4396] = -13'b0000010000100; // -132 -0.03216126188635826
storage[4397] = -13'b0000000000101; // -5 -0.001207191962748766
storage[4398] =  13'b0000000010011; // 19 0.004645434208214283
storage[4399] =  13'b0000010000111; // 135 0.03294771537184715
storage[4400] =  13'b0000001110000; // 112 0.02723539248108864
storage[4401] = -13'b0000001100100; // -100 -0.02448982372879982
storage[4402] =  13'b0000010101101; // 173 0.04233013466000557
storage[4403] = -13'b0000110111111; // -447 -0.10911483317613602
storage[4404] = -13'b0000000010111; // -23 -0.005628697108477354
storage[4405] = -13'b0000110110110; // -438 -0.1069808378815651
storage[4406] = -13'b0000001010000; // -80 -0.019478896632790565
storage[4407] =  13'b0000000011100; // 28 0.006950985640287399
storage[4408] =  13'b0000001101010; // 106 0.025973062962293625
storage[4409] =  13'b0000101010100; // 340 0.08309803903102875
storage[4410] =  13'b0000010010000; // 144 0.035130955278873444
storage[4411] =  13'b0000000111110; // 62 0.015086381696164608
storage[4412] =  13'b0000000101110; // 46 0.011197495274245739
storage[4413] =  13'b0000101011100; // 348 0.08498778194189072
storage[4414] =  13'b0000100001111; // 271 0.06606762111186981
storage[4415] = -13'b0000101011011; // -347 -0.08471405506134033
storage[4416] =  13'b0000110101100; // 428 0.10449793934822083
storage[4417] =  13'b0000001101100; // 108 0.026357604190707207
storage[4418] =  13'b0000011001010; // 202 0.049345798790454865
storage[4419] = -13'b0000000010000; // -16 -0.0040079141035676
storage[4420] = -13'b0001000001001; // -521 -0.12711940705776215
storage[4421] =  13'b0000000011000; // 24 0.0059132082387804985
storage[4422] = -13'b0000001010000; // -80 -0.019444629549980164
storage[4423] = -13'b0001100001000; // -776 -0.18950828909873962
storage[4424] = -13'b0001000111001; // -569 -0.13888481259346008
storage[4425] = -13'b0000110101101; // -429 -0.10463804751634598
storage[4426] = -13'b0000010111111; // -191 -0.04655035585165024
storage[4427] = -13'b0000110001111; // -399 -0.0973593071103096
storage[4428] = -13'b0000010100010; // -162 -0.039634186774492264
storage[4429] =  13'b0000100011100; // 284 0.06932241469621658
storage[4430] = -13'b0000000110100; // -52 -0.01264482643455267
storage[4431] = -13'b0000001011110; // -94 -0.02294214628636837
storage[4432] = -13'b0000010100101; // -165 -0.040383294224739075
storage[4433] =  13'b0000011101101; // 237 0.05790761113166809
storage[4434] =  13'b0000100010001; // 273 0.06662140041589737
storage[4435] =  13'b0000010011000; // 152 0.03701397404074669
storage[4436] = -13'b0000010100110; // -166 -0.040528565645217896
storage[4437] = -13'b0001011110111; // -759 -0.1853928416967392
storage[4438] =  13'b0000000011011; // 27 0.006547822616994381
storage[4439] =  13'b0000100010100; // 276 0.06736646592617035
storage[4440] = -13'b0000001100101; // -101 -0.024588337168097496
storage[4441] = -13'b0000000000100; // -4 -0.0008790249121375382
storage[4442] = -13'b0000010001001; // -137 -0.033373307436704636
storage[4443] =  13'b0000101101110; // 366 0.08928881585597992
storage[4444] =  13'b0000000100111; // 39 0.009417740628123283
storage[4445] = -13'b0000110010110; // -406 -0.0990893542766571
storage[4446] = -13'b0000011010100; // -212 -0.05173546075820923
storage[4447] =  13'b0000011001100; // 204 0.04980068281292915
storage[4448] = -13'b0000110111100; // -444 -0.10835745930671692
storage[4449] = -13'b0000000001010; // -10 -0.002548029413446784
storage[4450] =  13'b0000100111010; // 314 0.07674872875213623
storage[4451] = -13'b0000000111111; // -63 -0.015295437537133694
storage[4452] =  13'b0000001100001; // 97 0.023696094751358032
storage[4453] =  13'b0000101100110; // 358 0.0874660387635231
storage[4454] =  13'b0000001101100; // 108 0.02626749314367771
storage[4455] = -13'b0000000101000; // -40 -0.009780480526387691
storage[4456] = -13'b0000100110100; // -308 -0.07517438381910324
storage[4457] = -13'b0010000010000; // -1040 -0.2539510428905487
storage[4458] = -13'b0000110000000; // -384 -0.09386520087718964
storage[4459] = -13'b0001000010011; // -531 -0.1296670138835907
storage[4460] = -13'b0001101010000; // -848 -0.20712630450725555
storage[4461] = -13'b0001000100111; // -551 -0.13463160395622253
storage[4462] = -13'b0000010110110; // -182 -0.044536542147397995
storage[4463] =  13'b0000101100010; // 354 0.08641942590475082
storage[4464] = -13'b0000011001111; // -207 -0.05061902850866318
storage[4465] =  13'b0000001111100; // 124 0.030219068750739098
storage[4466] =  13'b0000011111101; // 253 0.06178756058216095
storage[4467] =  13'b0001000110101; // 565 0.13791148364543915
storage[4468] =  13'b0000000101000; // 40 0.009786047972738743
storage[4469] = -13'b0000001100000; // -96 -0.023483557626605034
storage[4470] =  13'b0001000010100; // 532 0.12994268536567688
storage[4471] =  13'b0000011110110; // 246 0.060097333043813705
storage[4472] = -13'b0000101000010; // -322 -0.07852014154195786
storage[4473] = -13'b0001010010001; // -657 -0.1603303700685501
storage[4474] = -13'b0000011000100; // -196 -0.04780391603708267
storage[4475] = -13'b0000001111001; // -121 -0.029566487297415733
storage[4476] =  13'b0000001000110; // 70 0.017108798027038574
storage[4477] = -13'b0000010000000; // -128 -0.031278081238269806
storage[4478] =  13'b0000000110000; // 48 0.011603853665292263
storage[4479] = -13'b0001011011010; // -730 -0.17811986804008484
storage[4480] = -13'b0001000100111; // -551 -0.1344357579946518
storage[4481] =  13'b0000010111010; // 186 0.04543834924697876
storage[4482] = -13'b0000100110001; // -305 -0.07441934943199158
storage[4483] =  13'b0000110001100; // 396 0.09675417840480804
storage[4484] =  13'b0000001100000; // 96 0.02341114729642868
storage[4485] = -13'b0001001001111; // -591 -0.14437972009181976
storage[4486] =  13'b0000100010111; // 279 0.06815649569034576
storage[4487] =  13'b0000010010001; // 145 0.03547092154622078
storage[4488] = -13'b0000111111110; // -510 -0.12452977150678635
storage[4489] = -13'b0000001110101; // -117 -0.028501244261860847
storage[4490] = -13'b0000110011010; // -410 -0.10002270340919495
storage[4491] = -13'b0000010101000; // -168 -0.04106675088405609
storage[4492] = -13'b0000100110101; // -309 -0.07550708204507828
storage[4493] = -13'b0000100110101; // -309 -0.07540279626846313
storage[4494] =  13'b0001010000001; // 641 0.15642023086547852
storage[4495] =  13'b0000011110110; // 246 0.05998745560646057
storage[4496] = -13'b0000001101100; // -108 -0.026261277496814728
storage[4497] =  13'b0000100010100; // 276 0.06745119392871857
storage[4498] = -13'b0000101101011; // -363 -0.08873408287763596
storage[4499] = -13'b0000100011111; // -287 -0.07001112401485443
storage[4500] = -13'b0001101101000; // -872 -0.21289537847042084
storage[4501] =  13'b0000010100100; // 164 0.03999597951769829
storage[4502] =  13'b0000000100111; // 39 0.009542935527861118
storage[4503] =  13'b0000010110000; // 176 0.04295250028371811
storage[4504] =  13'b0000011000100; // 196 0.04785388708114624
storage[4505] =  13'b0000001001111; // 79 0.019273728132247925
storage[4506] =  13'b0000101000101; // 325 0.07938408851623535
storage[4507] = -13'b0000001001010; // -74 -0.01812738925218582
storage[4508] = -13'b0000100111101; // -317 -0.07736096531152725
storage[4509] =  13'b0000111010000; // 464 0.11331748217344284
storage[4510] = -13'b0000010110000; // -176 -0.04305850714445114
storage[4511] = -13'b0000001001110; // -78 -0.018935516476631165
storage[4512] = -13'b0000011100000; // -224 -0.05470766872167587
storage[4513] =  13'b0000000101111; // 47 0.011544880457222462
storage[4514] =  13'b0000010000111; // 135 0.03302868828177452
storage[4515] =  13'b0000011110011; // 243 0.059295400977134705
storage[4516] =  13'b0000100100011; // 291 0.07115323096513748
storage[4517] =  13'b0000101000110; // 326 0.079536072909832
storage[4518] =  13'b0000001000100; // 68 0.016630161553621292
storage[4519] =  13'b0000111000001; // 449 0.10964952409267426
storage[4520] = -13'b0000100100010; // -290 -0.07078459858894348
storage[4521] = -13'b0000111001100; // -460 -0.11241301149129868
storage[4522] = -13'b0000011101000; // -232 -0.05666603147983551
storage[4523] = -13'b0000011111100; // -252 -0.06163962557911873
storage[4524] = -13'b0000001011010; // -90 -0.021959150210022926
storage[4525] = -13'b0000100110001; // -305 -0.07446711510419846
storage[4526] = -13'b0000011010100; // -212 -0.051771070808172226
storage[4527] = -13'b0000001011000; // -88 -0.021429764106869698
storage[4528] =  13'b0000110000111; // 391 0.09536553174257278
storage[4529] =  13'b0000100011100; // 284 0.06933658570051193
storage[4530] =  13'b0000001010110; // 86 0.02089023031294346
storage[4531] =  13'b0000101111000; // 376 0.09178676456212997
storage[4532] = -13'b0000011100110; // -230 -0.056030530482530594
storage[4533] = -13'b0000000011100; // -28 -0.006732504814863205
storage[4534] = -13'b0001001111010; // -634 -0.1547423005104065
storage[4535] = -13'b0001000100010; // -546 -0.13322196900844574
storage[4536] = -13'b0000110010100; // -404 -0.0986071303486824
storage[4537] =  13'b0000100100010; // 290 0.07083629816770554
storage[4538] = -13'b0000001101101; // -109 -0.026686623692512512
storage[4539] = -13'b0000011111011; // -251 -0.06123810634016991
storage[4540] =  13'b0000001010100; // 84 0.020400134846568108
storage[4541] =  13'b0000000110000; // 48 0.011828720569610596
storage[4542] = -13'b0000001010010; // -82 -0.02004271186888218
storage[4543] = -13'b0000101111010; // -378 -0.09236332029104233
storage[4544] =  13'b0000000111101; // 61 0.014922229573130608
storage[4545] =  13'b0000000111110; // 62 0.015096390619874
storage[4546] =  13'b0000111000100; // 452 0.11044865846633911
storage[4547] =  13'b0001001010111; // 599 0.1463385969400406
storage[4548] =  13'b0000011011110; // 222 0.05409757047891617
storage[4549] = -13'b0000010011111; // -159 -0.03872837498784065
storage[4550] =  13'b0000010001111; // 143 0.03482130914926529
storage[4551] = -13'b0000011011000; // -216 -0.05275159329175949
storage[4552] = -13'b0000011110010; // -242 -0.059123843908309937
storage[4553] = -13'b0001000011011; // -539 -0.13150528073310852
storage[4554] = -13'b0001001010001; // -593 -0.1448621153831482
storage[4555] = -13'b0000100011011; // -283 -0.0691993236541748
storage[4556] =  13'b0000001101010; // 106 0.025920487940311432
storage[4557] = -13'b0000110110111; // -439 -0.10714586824178696
storage[4558] = -13'b0000101010011; // -339 -0.08272972702980042
storage[4559] = -13'b0000101101110; // -366 -0.08942986279726028
storage[4560] = -13'b0000000000000; // 0 -4.791032915818505e-05
storage[4561] =  13'b0000011000100; // 196 0.04780271649360657
storage[4562] =  13'b0000010100101; // 165 0.04030745103955269
storage[4563] =  13'b0000110001011; // 395 0.09645276516675949
storage[4564] = -13'b0001100000111; // -775 -0.18918025493621826
storage[4565] =  13'b0000110000101; // 389 0.09487670660018921
storage[4566] =  13'b0000111101100; // 492 0.12023864686489105
storage[4567] = -13'b0001101100011; // -867 -0.2117205262184143
storage[4568] = -13'b0000101000011; // -323 -0.07875925302505493
storage[4569] =  13'b0000100010001; // 273 0.06654678285121918
storage[4570] = -13'b0001100000100; // -772 -0.18843452632427216
storage[4571] = -13'b0000010010001; // -145 -0.035457782447338104
storage[4572] = -13'b0000000001100; // -12 -0.002809748752042651
storage[4573] =  13'b0000011010100; // 212 0.051800038665533066
storage[4574] =  13'b0000010001000; // 136 0.033283915370702744
storage[4575] = -13'b0000110010011; // -403 -0.09832017123699188
storage[4576] =  13'b0000111100001; // 481 0.11742708086967468
storage[4577] =  13'b0001010011101; // 669 0.16339148581027985
storage[4578] = -13'b0010100001000; // -1288 -0.3143766522407532
storage[4579] = -13'b0000000000001; // -1 -0.0002212475228589028
storage[4580] = -13'b0000011100001; // -225 -0.05484020709991455
storage[4581] = -13'b0001101000110; // -838 -0.2046479433774948
storage[4582] =  13'b0000010001010; // 138 0.033733122050762177
storage[4583] =  13'b0000000001100; // 12 0.0029269265942275524
storage[4584] = -13'b0001000011110; // -542 -0.13230925798416138
storage[4585] =  13'b0000011101001; // 233 0.056917015463113785
storage[4586] =  13'b0000011110111; // 247 0.06025216355919838
storage[4587] = -13'b0000011111000; // -248 -0.06043723598122597
storage[4588] =  13'b0000000101101; // 45 0.010928056202828884
storage[4589] =  13'b0000000101101; // 45 0.010881147347390652
storage[4590] = -13'b0000110001101; // -397 -0.0968615934252739
storage[4591] = -13'b0000000011000; // -24 -0.005911475047469139
storage[4592] =  13'b0000111001101; // 461 0.11262129992246628
storage[4593] =  13'b0000001111001; // 121 0.02952505089342594
storage[4594] = -13'b0001110100111; // -935 -0.22838333249092102
storage[4595] = -13'b0001101110011; // -883 -0.21548601984977722
storage[4596] = -13'b0000100100011; // -291 -0.07103917747735977
storage[4597] = -13'b0000100001110; // -270 -0.06588000804185867
storage[4598] =  13'b0000000000001; // 1 0.0002969618944916874
storage[4599] =  13'b0000000000001; // 1 0.00012443576997611672
storage[4600] = -13'b0000000011100; // -28 -0.006766431964933872
storage[4601] =  13'b0000000101110; // 46 0.011203712783753872
storage[4602] = -13'b0000010010010; // -146 -0.03552637994289398
storage[4603] = -13'b0000101100110; // -358 -0.08732568472623825
storage[4604] = -13'b0001000100001; // -545 -0.13296134769916534
storage[4605] = -13'b0001011101011; // -747 -0.18242581188678741
storage[4606] = -13'b0000110101011; // -427 -0.10425137728452682
storage[4607] = -13'b0001000010111; // -535 -0.13051822781562805
storage[4608] =  13'b0000000110100; // 52 0.012792562134563923
storage[4609] =  13'b0000011010110; // 214 0.05216478556394577
storage[4610] =  13'b0000100110010; // 306 0.07471197098493576
storage[4611] = -13'b0000001010010; // -82 -0.020008902996778488
storage[4612] =  13'b0000011100101; // 229 0.05583664029836655
storage[4613] =  13'b0000010001101; // 141 0.03433912992477417
storage[4614] =  13'b0000110100001; // 417 0.10183484852313995
storage[4615] =  13'b0000001111111; // 127 0.030909841880202293
storage[4616] = -13'b0000010101011; // -171 -0.04176541790366173
storage[4617] =  13'b0000000000100; // 4 0.0010895599843934178
storage[4618] = -13'b0000101110010; // -370 -0.09040489792823792
storage[4619] = -13'b0001001110101; // -629 -0.1535748690366745
storage[4620] = -13'b0000110101000; // -424 -0.10357410460710526
storage[4621] = -13'b0001100101010; // -810 -0.19776834547519684
storage[4622] =  13'b0000000110000; // 48 0.011690392158925533
storage[4623] = -13'b0000001010101; // -85 -0.020632673054933548
storage[4624] = -13'b0001111111010; // -1018 -0.2485603541135788
storage[4625] = -13'b0000101110000; // -368 -0.08984265476465225
storage[4626] = -13'b0000010110001; // -177 -0.04322434216737747
storage[4627] = -13'b0000000111110; // -62 -0.01509476825594902
storage[4628] = -13'b0000000011010; // -26 -0.006423180922865868
storage[4629] = -13'b0000000110110; // -54 -0.013195772655308247
storage[4630] =  13'b0000001111110; // 126 0.030773665755987167
storage[4631] =  13'b0000110101010; // 426 0.10394430160522461
storage[4632] = -13'b0001001110011; // -627 -0.15308214724063873
storage[4633] = -13'b0000001101110; // -110 -0.026734573766589165
storage[4634] = -13'b0000000001010; // -10 -0.002513294806703925
storage[4635] = -13'b0010100111111; // -1343 -0.32797953486442566
storage[4636] =  13'b0000001110101; // 117 0.028567751869559288
storage[4637] = -13'b0000001110100; // -116 -0.028421126306056976
storage[4638] =  13'b0000010111000; // 184 0.0448274165391922
storage[4639] = -13'b0000000000111; // -7 -0.0016675599617883563
storage[4640] =  13'b0000000001010; // 10 0.0023425144609063864
storage[4641] = -13'b0010100100101; // -1317 -0.3214675784111023
storage[4642] = -13'b0000100101110; // -302 -0.07378311455249786
storage[4643] = -13'b0001111001101; // -973 -0.2376551777124405
storage[4644] = -13'b0001010110110; // -694 -0.1694549024105072
storage[4645] =  13'b0000001110100; // 116 0.028327133506536484
storage[4646] =  13'b0000001001000; // 72 0.01761518605053425
storage[4647] = -13'b0000000011000; // -24 -0.005938774440437555
storage[4648] =  13'b0000001111110; // 126 0.03078257292509079
storage[4649] =  13'b0000001010010; // 82 0.020042112097144127
storage[4650] =  13'b0000000101110; // 46 0.011233231984078884
storage[4651] =  13'b0000011111111; // 255 0.06220070645213127
storage[4652] = -13'b0000000000111; // -7 -0.0016400915337726474
storage[4653] = -13'b0010010011001; // -1177 -0.28736555576324463
storage[4654] =  13'b0000000000001; // 1 0.00022966056712903082
storage[4655] =  13'b0000010111011; // 187 0.0456385537981987
storage[4656] = -13'b0000011100101; // -229 -0.0557919479906559
storage[4657] =  13'b0000001011110; // 94 0.02299622632563114
storage[4658] =  13'b0000101100110; // 358 0.08749459683895111
storage[4659] = -13'b0000010111101; // -189 -0.04624726250767708
storage[4660] =  13'b0000010010010; // 146 0.03572635352611542
storage[4661] = -13'b0000101000010; // -322 -0.07849311083555222
storage[4662] = -13'b0000111111100; // -508 -0.12412156164646149
storage[4663] =  13'b0000000101100; // 44 0.010715053416788578
storage[4664] =  13'b0000001110110; // 118 0.028842555359005928
storage[4665] = -13'b0000010101010; // -170 -0.04143333062529564
storage[4666] =  13'b0001000010110; // 534 0.13026683032512665
storage[4667] =  13'b0000000111001; // 57 0.013857477344572544
storage[4668] = -13'b0001101010111; // -855 -0.20882068574428558
storage[4669] = -13'b0000101101101; // -365 -0.08903440088033676
storage[4670] =  13'b0000001111000; // 120 0.02932640351355076
storage[4671] =  13'b0000110001100; // 396 0.09661596268415451
storage[4672] =  13'b0000010110111; // 183 0.04456309229135513
storage[4673] =  13'b0000001011101; // 93 0.022667894139885902
storage[4674] =  13'b0000110011010; // 410 0.10011537373065948
storage[4675] =  13'b0000000111111; // 63 0.015261210501194
storage[4676] = -13'b0000011100111; // -231 -0.05631840229034424
storage[4677] = -13'b0001001110101; // -629 -0.15355601906776428
storage[4678] = -13'b0010010000110; // -1158 -0.2827225625514984
storage[4679] = -13'b0001010111101; // -701 -0.17104844748973846
storage[4680] = -13'b0001011011100; // -732 -0.17866021394729614
storage[4681] = -13'b0000000010110; // -22 -0.005362710449844599
storage[4682] =  13'b0000001000000; // 64 0.01572604849934578
storage[4683] =  13'b0000110110101; // 437 0.10663176327943802
storage[4684] = -13'b0000011100100; // -228 -0.055718425661325455
storage[4685] =  13'b0000001111110; // 126 0.030705949291586876
storage[4686] =  13'b0000011110100; // 244 0.05962860584259033
storage[4687] = -13'b0001111101100; // -1004 -0.24517884850502014
storage[4688] = -13'b0001110010001; // -913 -0.22291895747184753
storage[4689] = -13'b0010011001100; // -1228 -0.29970961809158325
storage[4690] = -13'b0000001011001; // -89 -0.021842459216713905
storage[4691] =  13'b0000001101000; // 104 0.025334177538752556
storage[4692] =  13'b0000110110011; // 435 0.10608100891113281
storage[4693] = -13'b0000010100000; // -160 -0.03909678012132645
storage[4694] = -13'b0000010101001; // -169 -0.04115027189254761
storage[4695] = -13'b0000101010001; // -337 -0.08216747641563416
storage[4696] = -13'b0000000001110; // -14 -0.0033714473247528076
storage[4697] = -13'b0000000010111; // -23 -0.005626797676086426
storage[4698] = -13'b0001100000101; // -773 -0.18879321217536926
storage[4699] =  13'b0000000000111; // 7 0.0017750808037817478
storage[4700] = -13'b0000001010100; // -84 -0.02049950137734413
storage[4701] = -13'b0000010001001; // -137 -0.03339337557554245
storage[4702] = -13'b0000000010111; // -23 -0.005534763913601637
storage[4703] =  13'b0000001000001; // 65 0.01586538925766945
storage[4704] = -13'b0000001000011; // -67 -0.016354458406567574
storage[4705] =  13'b0000100001000; // 264 0.06445103138685226
storage[4706] =  13'b0000010100100; // 164 0.04002753645181656
storage[4707] = -13'b0000011110011; // -243 -0.059287384152412415
storage[4708] = -13'b0000100001011; // -267 -0.06522119045257568
storage[4709] = -13'b0000101111000; // -376 -0.09178618341684341
storage[4710] =  13'b0000000010010; // 18 0.004361523315310478
storage[4711] = -13'b0000001110011; // -115 -0.0279629398137331
storage[4712] = -13'b0000110111110; // -446 -0.10890676826238632
storage[4713] = -13'b0000111101000; // -488 -0.119180828332901
storage[4714] = -13'b0000010000010; // -130 -0.03179318457841873
storage[4715] = -13'b0000100111011; // -315 -0.07695192843675613
storage[4716] =  13'b0000000000010; // 2 0.0004753510293085128
storage[4717] = -13'b0000001111000; // -120 -0.029373381286859512
storage[4718] = -13'b0000000101010; // -42 -0.010302855633199215
storage[4719] = -13'b0000010110001; // -177 -0.04311829432845116
storage[4720] =  13'b0000011000111; // 199 0.04856691136956215
storage[4721] =  13'b0000000010010; // 18 0.004432643763720989
storage[4722] =  13'b0000000101001; // 41 0.010081361047923565
storage[4723] = -13'b0000111001101; // -461 -0.112607941031456
storage[4724] =  13'b0000101100100; // 356 0.08693088591098785
storage[4725] = -13'b0000010111111; // -191 -0.04661446809768677
storage[4726] = -13'b0000011010100; // -212 -0.05179004743695259
storage[4727] = -13'b0000001010001; // -81 -0.019709469750523567
storage[4728] = -13'b0000011001011; // -203 -0.04945674538612366
storage[4729] = -13'b0000000100101; // -37 -0.009001458995044231
storage[4730] =  13'b0000100110000; // 304 0.07418831437826157
storage[4731] =  13'b0000010010010; // 146 0.03563375771045685
storage[4732] =  13'b0000001001001; // 73 0.01771102473139763
storage[4733] =  13'b0000011011010; // 218 0.05312759801745415
storage[4734] = -13'b0000010110000; // -176 -0.04302358627319336
storage[4735] = -13'b0001000000110; // -518 -0.12646692991256714
storage[4736] = -13'b0001000100000; // -544 -0.13271136581897736
storage[4737] = -13'b0000100100000; // -288 -0.0703861340880394
storage[4738] = -13'b0010000001001; // -1033 -0.2520880401134491
storage[4739] = -13'b0001010110011; // -691 -0.1687716394662857
storage[4740] = -13'b0000011010111; // -215 -0.05251792445778847
storage[4741] = -13'b0000110011000; // -408 -0.09963558614253998
storage[4742] =  13'b0000001101111; // 111 0.027132075279951096
storage[4743] =  13'b0000000001001; // 9 0.0022567673586308956
storage[4744] =  13'b0000100001111; // 271 0.06609419733285904
storage[4745] =  13'b0000000111110; // 62 0.015204491093754768
storage[4746] = -13'b0000110001111; // -399 -0.09734214097261429
storage[4747] = -13'b0000000000000; // 0 -0.00011234464182052761
storage[4748] = -13'b0000010010110; // -150 -0.03670595958828926
storage[4749] = -13'b0001000100101; // -549 -0.13397498428821564
storage[4750] = -13'b0000010101011; // -171 -0.041646674275398254
storage[4751] = -13'b0000010101010; // -170 -0.04152694717049599
storage[4752] =  13'b0000010100010; // 162 0.03961985185742378
storage[4753] = -13'b0000001010001; // -81 -0.019753871485590935
storage[4754] =  13'b0000100100100; // 292 0.07140941917896271
storage[4755] =  13'b0000100011011; // 283 0.06916457414627075
storage[4756] =  13'b0000000100011; // 35 0.008445460349321365
storage[4757] = -13'b0000000110110; // -54 -0.013302060775458813
storage[4758] =  13'b0000100010010; // 274 0.06688534468412399
storage[4759] =  13'b0000101000101; // 325 0.07945965975522995
storage[4760] = -13'b0000001000101; // -69 -0.01679920218884945
storage[4761] = -13'b0000000000110; // -6 -0.0013821288011968136
storage[4762] =  13'b0000111100110; // 486 0.11876554787158966
storage[4763] =  13'b0000011101101; // 237 0.057824768126010895
storage[4764] =  13'b0000111111000; // 504 0.12293842434883118
storage[4765] =  13'b0000000111101; // 61 0.014955724589526653
storage[4766] = -13'b0000010011110; // -158 -0.03850643336772919
storage[4767] = -13'b0000100101000; // -296 -0.0722164735198021
storage[4768] =  13'b0000101001101; // 333 0.08132883906364441
storage[4769] = -13'b0000010101101; // -173 -0.042352475225925446
storage[4770] = -13'b0000010000001; // -129 -0.031419672071933746
storage[4771] = -13'b0000010000100; // -132 -0.032206472009420395
storage[4772] =  13'b0000010101010; // 170 0.041414931416511536
storage[4773] =  13'b0000011110001; // 241 0.05876987800002098
storage[4774] =  13'b0000011110101; // 245 0.059738077223300934
storage[4775] =  13'b0000101010010; // 338 0.08248468488454819
storage[4776] =  13'b0000010111010; // 186 0.04549175500869751
storage[4777] =  13'b0000100100010; // 290 0.07076333463191986
storage[4778] =  13'b0000100010100; // 276 0.06734804064035416
storage[4779] =  13'b0000010001011; // 139 0.03391711413860321
storage[4780] =  13'b0001001101010; // 618 0.15096507966518402
storage[4781] =  13'b0000010001111; // 143 0.03482942655682564
storage[4782] =  13'b0000000010111; // 23 0.005680386908352375
storage[4783] =  13'b0000001011101; // 93 0.022790955379605293
storage[4784] = -13'b0000101010000; // -336 -0.08213900774717331
storage[4785] =  13'b0000001100010; // 98 0.023855509236454964
storage[4786] =  13'b0000101001010; // 330 0.08045055717229843
storage[4787] = -13'b0000011000111; // -199 -0.0485982708632946
storage[4788] =  13'b0000101100100; // 356 0.086935855448246
storage[4789] = -13'b0010000111111; // -1087 -0.2653033435344696
storage[4790] = -13'b0010011011011; // -1243 -0.3035130202770233
storage[4791] = -13'b0001000000100; // -516 -0.12607327103614807
storage[4792] =  13'b0001000110001; // 561 0.13698551058769226
storage[4793] = -13'b0000001100110; // -102 -0.024934949353337288
storage[4794] =  13'b0000100101000; // 296 0.07228588312864304
storage[4795] =  13'b0001000011011; // 539 0.13159707188606262
storage[4796] =  13'b0000110100001; // 417 0.1019132062792778
storage[4797] =  13'b0000100110001; // 305 0.07442952692508698
storage[4798] = -13'b0000101000111; // -327 -0.07983507961034775
storage[4799] = -13'b0001000101100; // -556 -0.13576751947402954
storage[4800] = -13'b0001101001111; // -847 -0.2068883776664734
storage[4801] =  13'b0000010001010; // 138 0.0335959829390049
storage[4802] = -13'b0000010101111; // -175 -0.0426938533782959
storage[4803] = -13'b0000111000000; // -448 -0.10946246236562729
storage[4804] =  13'b0000011010100; // 212 0.05166172608733177
storage[4805] =  13'b0000010010111; // 151 0.0369587242603302
storage[4806] =  13'b0000001100011; // 99 0.02424255572259426
storage[4807] = -13'b0000100001111; // -271 -0.06612187623977661
storage[4808] = -13'b0000000100000; // -32 -0.007880003191530704
storage[4809] = -13'b0000000011000; // -24 -0.005900188814848661
storage[4810] = -13'b0000000110101; // -53 -0.013058231212198734
storage[4811] =  13'b0000101011001; // 345 0.08413547277450562
storage[4812] = -13'b0000000000011; // -3 -0.0006456763367168605
storage[4813] = -13'b0000010111010; // -186 -0.04529160261154175
storage[4814] =  13'b0000001100000; // 96 0.02351919375360012
storage[4815] =  13'b0000100100101; // 293 0.07161150127649307
storage[4816] =  13'b0000010001011; // 139 0.0338745079934597
storage[4817] = -13'b0000001001010; // -74 -0.018100328743457794
storage[4818] = -13'b0000010111010; // -186 -0.04546486586332321
storage[4819] =  13'b0000000101100; // 44 0.010684769600629807
storage[4820] = -13'b0000000101000; // -40 -0.009836276061832905
storage[4821] = -13'b0000000110000; // -48 -0.011677426286041737
storage[4822] =  13'b0000100011110; // 286 0.06988371163606644
storage[4823] =  13'b0000011010110; // 214 0.052193716168403625
storage[4824] = -13'b0000011001111; // -207 -0.05062951147556305
storage[4825] =  13'b0000001001111; // 79 0.019266366958618164
storage[4826] = -13'b0000101010111; // -343 -0.08366712927818298
storage[4827] = -13'b0000010010111; // -151 -0.03696691244840622
storage[4828] =  13'b0000010110110; // 182 0.04431269317865372
storage[4829] =  13'b0000000001000; // 8 0.00207171100191772
storage[4830] =  13'b0000000101011; // 43 0.010388748720288277
storage[4831] =  13'b0000111101111; // 495 0.12078433483839035
storage[4832] = -13'b0000001100100; // -100 -0.02436145953834057
storage[4833] = -13'b0000001100101; // -101 -0.02459901012480259
storage[4834] = -13'b0000010010000; // -144 -0.03520715609192848
storage[4835] = -13'b0000110010000; // -400 -0.09754263609647751
storage[4836] = -13'b0010000101101; // -1069 -0.26096025109291077
storage[4837] = -13'b0000000010000; // -16 -0.003853857982903719
storage[4838] = -13'b0000100010001; // -273 -0.06669443845748901
storage[4839] = -13'b0001000010100; // -532 -0.12983570992946625
storage[4840] =  13'b0000011101110; // 238 0.058033913373947144
storage[4841] =  13'b0000001110110; // 118 0.028920114040374756
storage[4842] = -13'b0000010101001; // -169 -0.041379135102033615
storage[4843] = -13'b0000111001011; // -459 -0.11213897168636322
storage[4844] = -13'b0000001100001; // -97 -0.02379530668258667
storage[4845] = -13'b0000111011110; // -478 -0.11661416292190552
storage[4846] = -13'b0001000100001; // -545 -0.13297507166862488
storage[4847] = -13'b0000100100001; // -289 -0.07051481306552887
storage[4848] = -13'b0001010000101; // -645 -0.15738064050674438
storage[4849] =  13'b0000000101110; // 46 0.011160075664520264
storage[4850] = -13'b0000000001111; // -15 -0.0036042651627212763
storage[4851] = -13'b0001001011111; // -607 -0.14826977252960205
storage[4852] = -13'b0000111110100; // -500 -0.12196488678455353
storage[4853] = -13'b0000100011111; // -287 -0.07003732770681381
storage[4854] = -13'b0000011011001; // -217 -0.05295857787132263
storage[4855] = -13'b0001000011001; // -537 -0.1311596781015396
storage[4856] =  13'b0000011001101; // 205 0.0499558262526989
storage[4857] =  13'b0000011010111; // 215 0.052369944751262665
storage[4858] = -13'b0000001111111; // -127 -0.030979618430137634
storage[4859] =  13'b0000100000001; // 257 0.06277173012495041
storage[4860] =  13'b0000101001010; // 330 0.08053640276193619
storage[4861] = -13'b0000010100010; // -162 -0.039609793573617935
storage[4862] = -13'b0000000000110; // -6 -0.0015826483722776175
storage[4863] =  13'b0000001111100; // 124 0.030302276834845543
storage[4864] =  13'b0000001110110; // 118 0.02876126579940319
storage[4865] =  13'b0000010001011; // 139 0.03388656675815582
storage[4866] =  13'b0000100101000; // 296 0.07215440273284912
storage[4867] =  13'b0000011001001; // 201 0.049157749861478806
storage[4868] =  13'b0000001010010; // 82 0.0199167188256979
storage[4869] =  13'b0000011010010; // 210 0.05118982493877411
storage[4870] =  13'b0000000110110; // 54 0.013188307173550129
storage[4871] =  13'b0000100010101; // 277 0.06763271242380142
storage[4872] =  13'b0000001000101; // 69 0.016768572852015495
storage[4873] =  13'b0000001100000; // 96 0.02333703264594078
storage[4874] = -13'b0000010100000; // -160 -0.0391518771648407
storage[4875] =  13'b0000101000011; // 323 0.0787639170885086
storage[4876] = -13'b0000010000110; // -134 -0.03261241316795349
storage[4877] = -13'b0000100001100; // -268 -0.06537413597106934
storage[4878] =  13'b0000010010001; // 145 0.03530662879347801
storage[4879] =  13'b0000000100100; // 36 0.008753218688070774
storage[4880] =  13'b0000100101011; // 299 0.07294926047325134
storage[4881] =  13'b0000011100001; // 225 0.054845843464136124
storage[4882] =  13'b0000101000110; // 326 0.07962549477815628
storage[4883] =  13'b0000100110011; // 307 0.07500553876161575
storage[4884] = -13'b0000001000110; // -70 -0.017172403633594513
storage[4885] = -13'b0001001001100; // -588 -0.1436314582824707
storage[4886] = -13'b0001110001101; // -909 -0.22190895676612854
storage[4887] = -13'b0000010100001; // -161 -0.039206065237522125
storage[4888] = -13'b0000000000001; // -1 -0.000311883952235803
storage[4889] = -13'b0000101100100; // -356 -0.0869329571723938
storage[4890] = -13'b0010001111111; // -1151 -0.2808944880962372
storage[4891] = -13'b0000011100101; // -229 -0.05581814795732498
storage[4892] = -13'b0000100010010; // -274 -0.06691437214612961
storage[4893] =  13'b0000011100110; // 230 0.05626223236322403
storage[4894] =  13'b0000001111111; // 127 0.0309771578758955
storage[4895] = -13'b0000000000001; // -1 -0.0002603247994557023
storage[4896] =  13'b0000110100100; // 420 0.10260093212127686
storage[4897] =  13'b0000001100110; // 102 0.024808932095766068
storage[4898] =  13'b0000010011101; // 157 0.03830885887145996
storage[4899] =  13'b0000101001101; // 333 0.08128035813570023
storage[4900] =  13'b0000101100001; // 353 0.08614695817232132
storage[4901] = -13'b0000100010010; // -274 -0.06684275716543198
storage[4902] = -13'b0000101101000; // -360 -0.08800148218870163
storage[4903] =  13'b0000010010110; // 150 0.03671514615416527
storage[4904] =  13'b0000010100101; // 165 0.04039692133665085
storage[4905] =  13'b0000011110001; // 241 0.05880706012248993
storage[4906] =  13'b0000001001110; // 78 0.019123660400509834
storage[4907] = -13'b0000011010011; // -211 -0.05153263732790947
storage[4908] = -13'b0000001001110; // -78 -0.01899447664618492
storage[4909] = -13'b0001111110101; // -1013 -0.24721233546733856
storage[4910] = -13'b0000100010011; // -275 -0.06718740612268448
storage[4911] = -13'b0000000111101; // -61 -0.014881000854074955
storage[4912] = -13'b0000011101110; // -238 -0.058213479816913605
storage[4913] =  13'b0000001111000; // 120 0.02920941449701786
storage[4914] = -13'b0000001100011; // -99 -0.024214597418904305
storage[4915] = -13'b0000000011101; // -29 -0.007094722241163254
storage[4916] = -13'b0000001101001; // -105 -0.025683648884296417
storage[4917] = -13'b0000000101111; // -47 -0.011510724201798439
storage[4918] = -13'b0000100010101; // -277 -0.06773427128791809
storage[4919] =  13'b0000010101010; // 170 0.041569165885448456
storage[4920] =  13'b0000010011011; // 155 0.0378534272313118
storage[4921] =  13'b0000101011000; // 344 0.08387890458106995
storage[4922] =  13'b0000011110001; // 241 0.05889159440994263
storage[4923] =  13'b0000011011001; // 217 0.05288053676486015
storage[4924] =  13'b0000000111100; // 60 0.014581575989723206
storage[4925] = -13'b0000001100101; // -101 -0.024633053690195084
storage[4926] = -13'b0000001000010; // -66 -0.01618254743516445
storage[4927] = -13'b0000111110100; // -500 -0.12213952839374542
storage[4928] = -13'b0001001010101; // -597 -0.14565598964691162
storage[4929] = -13'b0000010010110; // -150 -0.03654598444700241
storage[4930] = -13'b0000001000000; // -64 -0.01554812677204609
storage[4931] = -13'b0000001010001; // -81 -0.01973886787891388
storage[4932] =  13'b0000110101001; // 425 0.10384413599967957
storage[4933] = -13'b0000000111111; // -63 -0.015468495897948742
storage[4934] = -13'b0000010001100; // -140 -0.03423476591706276
storage[4935] = -13'b0000000001100; // -12 -0.0028493523132056
storage[4936] = -13'b0000001010010; // -82 -0.020119646564126015
storage[4937] = -13'b0001001101111; // -623 -0.152115136384964
storage[4938] =  13'b0000011011111; // 223 0.05451434478163719
storage[4939] = -13'b0000111101000; // -488 -0.11924371123313904
storage[4940] = -13'b0000111100011; // -483 -0.1178579032421112
storage[4941] =  13'b0000010010000; // 144 0.035090889781713486
storage[4942] = -13'b0000001100000; // -96 -0.0234361719340086
storage[4943] =  13'b0000100011001; // 281 0.06855334341526031
storage[4944] =  13'b0001000011001; // 537 0.1312035769224167
storage[4945] = -13'b0000000110110; // -54 -0.013277443125844002
storage[4946] =  13'b0000000111111; // 63 0.015500275418162346
storage[4947] =  13'b0000100001100; // 268 0.0654781311750412
storage[4948] = -13'b0000101111101; // -381 -0.09298989176750183
storage[4949] = -13'b0000011010110; // -214 -0.05236752703785896
storage[4950] = -13'b0000011110100; // -244 -0.05960437282919884
storage[4951] = -13'b0000011111111; // -255 -0.062149226665496826
storage[4952] =  13'b0000001011110; // 94 0.022916797548532486
storage[4953] =  13'b0000011100000; // 224 0.05477611720561981
storage[4954] =  13'b0000001010111; // 87 0.02112990990281105
storage[4955] = -13'b0000001010000; // -80 -0.019649198278784752
storage[4956] = -13'b0001010100001; // -673 -0.16422909498214722
storage[4957] =  13'b0001000101100; // 556 0.13566987216472626
storage[4958] =  13'b0000100110101; // 309 0.07546403259038925
storage[4959] =  13'b0000010100111; // 167 0.04087947681546211
storage[4960] =  13'b0000111000011; // 451 0.11015036702156067
storage[4961] =  13'b0000010000000; // 128 0.03126397356390953
storage[4962] = -13'b0000000001100; // -12 -0.002831675810739398
storage[4963] = -13'b0001011000111; // -711 -0.17347466945648193
storage[4964] =  13'b0000000100100; // 36 0.008830154314637184
storage[4965] =  13'b0000001110000; // 112 0.0273931585252285
storage[4966] = -13'b0001010001100; // -652 -0.1592697650194168
storage[4967] = -13'b0000010100001; // -161 -0.03927664831280708
storage[4968] =  13'b0000001011110; // 94 0.023052167147397995
storage[4969] =  13'b0000100111011; // 315 0.07683414965867996
storage[4970] = -13'b0000010010111; // -151 -0.03692205250263214
storage[4971] =  13'b0000101100111; // 359 0.08766775578260422
storage[4972] = -13'b0001101010101; // -853 -0.20831432938575745
storage[4973] = -13'b0000001010011; // -83 -0.0202837735414505
storage[4974] =  13'b0001000110101; // 565 0.13782216608524323
storage[4975] = -13'b0001000000110; // -518 -0.12655985355377197
storage[4976] =  13'b0000110011111; // 415 0.10129373520612717
storage[4977] =  13'b0000011110011; // 243 0.05924254655838013
storage[4978] = -13'b0000001110000; // -112 -0.02734196186065674
storage[4979] =  13'b0000001000000; // 64 0.015615592710673809
storage[4980] =  13'b0000101100010; // 354 0.08643560856580734
storage[4981] =  13'b0000011110101; // 245 0.05974884703755379
storage[4982] =  13'b0000100010110; // 278 0.0678640678524971
storage[4983] =  13'b0000100011000; // 280 0.06826967746019363
storage[4984] = -13'b0000100010101; // -277 -0.06771500408649445
storage[4985] = -13'b0000100001110; // -270 -0.0659153088927269
storage[4986] = -13'b0000001101010; // -106 -0.025979021564126015
storage[4987] = -13'b0000000100010; // -34 -0.008283279836177826
storage[4988] = -13'b0000001101000; // -104 -0.02531363256275654
storage[4989] = -13'b0000101110110; // -374 -0.091342031955719
storage[4990] =  13'b0000110010100; // 404 0.09861671179533005
storage[4991] =  13'b0000110110010; // 434 0.1058763638138771
storage[4992] = -13'b0000001000011; // -67 -0.01643221080303192
storage[4993] =  13'b0000000011001; // 25 0.006050820462405682
storage[4994] = -13'b0000100101111; // -303 -0.07396681606769562
storage[4995] = -13'b0001001000101; // -581 -0.1419123113155365
storage[4996] = -13'b0000000101110; // -46 -0.011275841854512691
storage[4997] =  13'b0000001011001; // 89 0.021841224282979965
storage[4998] =  13'b0000010101110; // 174 0.04254624620079994
storage[4999] = -13'b0000001000001; // -65 -0.01574805937707424
storage[5000] = -13'b0000010111000; // -184 -0.04492335394024849
storage[5001] =  13'b0000001001010; // 74 0.018017539754509926
storage[5002] = -13'b0000111101111; // -495 -0.12075802683830261
storage[5003] = -13'b0001001100100; // -612 -0.14942413568496704
storage[5004] = -13'b0000101111110; // -382 -0.09334476292133331
storage[5005] =  13'b0000011101100; // 236 0.0576254203915596
storage[5006] = -13'b0000101011111; // -351 -0.0857560858130455
storage[5007] = -13'b0010001001001; // -1097 -0.2677399218082428
storage[5008] = -13'b0001110001100; // -908 -0.22156037390232086
storage[5009] = -13'b0000011111101; // -253 -0.06168482452630997
storage[5010] = -13'b0000101001101; // -333 -0.08118699491024017
storage[5011] = -13'b0001101100011; // -867 -0.21158893406391144
storage[5012] = -13'b0001111000001; // -961 -0.23462210595607758
storage[5013] =  13'b0000000110110; // 54 0.013145465403795242
storage[5014] =  13'b0000001110010; // 114 0.027787717059254646
storage[5015] =  13'b0000010001010; // 138 0.033620234578847885
storage[5016] = -13'b0000110100011; // -419 -0.1021895632147789
storage[5017] =  13'b0000100001001; // 265 0.06476397067308426
storage[5018] =  13'b0000000010110; // 22 0.005409564822912216
storage[5019] = -13'b0001100000010; // -770 -0.187929168343544
storage[5020] = -13'b0000110100010; // -418 -0.10193156450986862
storage[5021] = -13'b0000110110101; // -437 -0.10660485923290253
storage[5022] =  13'b0000001011010; // 90 0.021974753588438034
storage[5023] = -13'b0000010101011; // -171 -0.041720885783433914
storage[5024] =  13'b0000011111101; // 253 0.061695653945207596
storage[5025] =  13'b0000011111100; // 252 0.06141161918640137
storage[5026] =  13'b0000001111101; // 125 0.030410774052143097
storage[5027] =  13'b0000100111000; // 312 0.07605382800102234
storage[5028] =  13'b0000001010110; // 86 0.020990123972296715
storage[5029] =  13'b0000001110111; // 119 0.029029754921793938
storage[5030] =  13'b0000000111111; // 63 0.015304045751690865
storage[5031] = -13'b0000101110000; // -368 -0.08974573016166687
storage[5032] =  13'b0000001101010; // 106 0.025843191891908646
storage[5033] = -13'b0001001100111; // -615 -0.15003973245620728
storage[5034] =  13'b0000101101100; // 364 0.08887002617120743
storage[5035] = -13'b0000001011111; // -95 -0.0232622642070055
storage[5036] = -13'b0000010000111; // -135 -0.032853689044713974
storage[5037] =  13'b0000111101010; // 490 0.11954020708799362
storage[5038] =  13'b0000111000100; // 452 0.11029694974422455
storage[5039] =  13'b0000111101110; // 494 0.1205231100320816
storage[5040] = -13'b0000000111010; // -58 -0.014132496900856495
storage[5041] =  13'b0001000100100; // 548 0.13370154798030853
storage[5042] =  13'b0000100100011; // 291 0.07101552933454514
storage[5043] = -13'b0000010111111; // -191 -0.04657869040966034
storage[5044] =  13'b0001010000110; // 646 0.1577494740486145
storage[5045] =  13'b0000011000100; // 196 0.04776538163423538
storage[5046] = -13'b0000000101110; // -46 -0.011160854250192642
storage[5047] = -13'b0001011001110; // -718 -0.17524240911006927
storage[5048] = -13'b0000010011000; // -152 -0.03704783320426941
storage[5049] =  13'b0000100110111; // 311 0.07591839879751205
storage[5050] = -13'b0000010001001; // -137 -0.033348433673381805
storage[5051] =  13'b0000011111010; // 250 0.061130769550800323
storage[5052] = -13'b0000111010110; // -470 -0.11466199159622192
storage[5053] =  13'b0000010011010; // 154 0.03765648975968361
storage[5054] = -13'b0000110011011; // -411 -0.10021989047527313
storage[5055] = -13'b0000010100100; // -164 -0.040123771876096725
storage[5056] = -13'b0000000010111; // -23 -0.005579962860792875
storage[5057] = -13'b0000011000111; // -199 -0.048499174416065216
storage[5058] = -13'b0001101010011; // -851 -0.20772798359394073
storage[5059] = -13'b0000011100100; // -228 -0.05557656288146973
storage[5060] = -13'b0001000101100; // -556 -0.13563528656959534
storage[5061] = -13'b0010011101100; // -1260 -0.3075914978981018
storage[5062] =  13'b0000001000001; // 65 0.015974976122379303
storage[5063] = -13'b0000110000101; // -389 -0.09489045292139053
storage[5064] = -13'b0001001000001; // -577 -0.14081740379333496
storage[5065] = -13'b0001000100110; // -550 -0.13428187370300293
storage[5066] = -13'b0000010001010; // -138 -0.0336422473192215
storage[5067] = -13'b0001011010011; // -723 -0.17643596231937408
storage[5068] =  13'b0001100110100; // 820 0.2002207338809967
storage[5069] = -13'b0000011010011; // -211 -0.05157534033060074
storage[5070] =  13'b0000101001011; // 331 0.08075104653835297
storage[5071] = -13'b0000111110001; // -497 -0.12134969979524612
storage[5072] = -13'b0001110100011; // -931 -0.22721149027347565
storage[5073] =  13'b0000001101010; // 106 0.02584490180015564
storage[5074] = -13'b0000010110000; // -176 -0.04304641857743263
storage[5075] =  13'b0000000110100; // 52 0.012711834162473679
storage[5076] = -13'b0000010010110; // -150 -0.036695171147584915
storage[5077] =  13'b0000000010111; // 23 0.005720375571399927
storage[5078] =  13'b0000100001100; // 268 0.06539689749479294
storage[5079] =  13'b0000000010001; // 17 0.004239865578711033
storage[5080] = -13'b0000001001110; // -78 -0.01900719664990902
storage[5081] = -13'b0000010111100; // -188 -0.04596089944243431
storage[5082] = -13'b0001000001101; // -525 -0.1282687932252884
storage[5083] = -13'b0001001010111; // -599 -0.14631043374538422
storage[5084] = -13'b0001011011010; // -730 -0.17826725542545319
storage[5085] = -13'b0000110010011; // -403 -0.09847262501716614
storage[5086] = -13'b0000000101110; // -46 -0.011198201216757298
storage[5087] = -13'b0000001000001; // -65 -0.015845833346247673
storage[5088] =  13'b0000001000000; // 64 0.015729518607258797
storage[5089] = -13'b0000001011011; // -91 -0.022188257426023483
storage[5090] =  13'b0000011011010; // 218 0.05322317034006119
storage[5091] = -13'b0000010001111; // -143 -0.03487459942698479
storage[5092] = -13'b0000000111010; // -58 -0.014122424647212029
storage[5093] = -13'b0000111001010; // -458 -0.11193311214447021
storage[5094] =  13'b0000000011111; // 31 0.007682671304792166
storage[5095] =  13'b0001000000111; // 519 0.1266784965991974
storage[5096] =  13'b0000011100000; // 224 0.05471761152148247
storage[5097] = -13'b0000011010111; // -215 -0.052444953471422195
storage[5098] =  13'b0000001111100; // 124 0.03025631420314312
storage[5099] = -13'b0001011011101; // -733 -0.17894048988819122
storage[5100] =  13'b0000101010011; // 339 0.08284229040145874
storage[5101] = -13'b0000110111110; // -446 -0.10878250747919083
storage[5102] =  13'b0000001110011; // 115 0.028119593858718872
storage[5103] = -13'b0000000100011; // -35 -0.008655337616801262
storage[5104] = -13'b0000011100010; // -226 -0.05519215390086174
storage[5105] = -13'b0000011010101; // -213 -0.05190061777830124
storage[5106] = -13'b0000011111101; // -253 -0.06171218678355217
storage[5107] = -13'b0000000010111; // -23 -0.005599382799118757
storage[5108] =  13'b0000000101000; // 40 0.009718412533402443
storage[5109] = -13'b0001110010000; // -912 -0.22260382771492004
storage[5110] = -13'b0001000101000; // -552 -0.13475361466407776
storage[5111] = -13'b0000111001000; // -456 -0.11129381507635117
storage[5112] = -13'b0001000101000; // -552 -0.13472288846969604
storage[5113] =  13'b0000010100001; // 161 0.039425864815711975
storage[5114] =  13'b0000001100011; // 99 0.02427954599261284
storage[5115] = -13'b0000101000110; // -326 -0.07958698272705078
storage[5116] =  13'b0000010010100; // 148 0.036226555705070496
storage[5117] = -13'b0000111111001; // -505 -0.12323478609323502
storage[5118] = -13'b0010010000110; // -1158 -0.2827768921852112
storage[5119] = -13'b0001001011001; // -601 -0.14662007987499237
storage[5120] = -13'b0010010100001; // -1185 -0.28930583596229553
storage[5121] = -13'b0001100010110; // -790 -0.1928885579109192
storage[5122] =  13'b0000110011110; // 414 0.10098965466022491
storage[5123] =  13'b0001001000100; // 580 0.14148133993148804
storage[5124] = -13'b0001100001011; // -779 -0.19007207453250885
storage[5125] = -13'b0000000010010; // -18 -0.004446758888661861
storage[5126] = -13'b0000100101010; // -298 -0.0727190151810646
storage[5127] = -13'b0010011110011; // -1267 -0.3092566430568695
storage[5128] =  13'b0000000000011; // 3 0.0007824643398635089
storage[5129] = -13'b0000110110110; // -438 -0.10685314983129501
storage[5130] = -13'b0000100010110; // -278 -0.0679522454738617
storage[5131] =  13'b0000001011010; // 90 0.022012602537870407
storage[5132] = -13'b0000010111011; // -187 -0.0457298718392849
storage[5133] = -13'b0000010100110; // -166 -0.0406075119972229
storage[5134] =  13'b0000001111011; // 123 0.029948066920042038
storage[5135] = -13'b0000110010111; // -407 -0.09930771589279175
storage[5136] = -13'b0000101101001; // -361 -0.08817650377750397
storage[5137] =  13'b0000000111001; // 57 0.014010350219905376
storage[5138] = -13'b0000101110001; // -369 -0.09011173248291016
storage[5139] = -13'b0000110010110; // -406 -0.09900271147489548
storage[5140] = -13'b0001010001100; // -652 -0.15915846824645996
storage[5141] = -13'b0000111110001; // -497 -0.1214008703827858
storage[5142] = -13'b0000011000011; // -195 -0.04755491018295288
storage[5143] = -13'b0000111001001; // -457 -0.11156461387872696
storage[5144] = -13'b0000100011100; // -284 -0.06944707781076431
storage[5145] =  13'b0000000010101; // 21 0.0052442243322730064
storage[5146] = -13'b0000001111110; // -126 -0.03075101226568222
storage[5147] =  13'b0000011100010; // 226 0.05509522929787636
storage[5148] =  13'b0000101100000; // 352 0.08584057539701462
storage[5149] = -13'b0000001110001; // -113 -0.027675101533532143
storage[5150] =  13'b0000101011000; // 344 0.08394481986761093
storage[5151] =  13'b0000011111111; // 255 0.06222367286682129
storage[5152] = -13'b0001100000101; // -773 -0.188822403550148
storage[5153] =  13'b0000000011110; // 30 0.007444930262863636
storage[5154] =  13'b0000010110001; // 177 0.04312998428940773
storage[5155] = -13'b0000100100001; // -289 -0.0705522894859314
storage[5156] =  13'b0000101001000; // 328 0.08003216981887817
storage[5157] =  13'b0000100000111; // 263 0.06414791196584702
storage[5158] =  13'b0000010111111; // 191 0.04655329883098602
storage[5159] = -13'b0000111000111; // -455 -0.11101806908845901
storage[5160] = -13'b0000111100110; // -486 -0.11858538538217545
storage[5161] = -13'b0000000001010; // -10 -0.002413193928077817
storage[5162] = -13'b0000000011111; // -31 -0.007460196502506733
storage[5163] = -13'b0000011100000; // -224 -0.05473996326327324
storage[5164] =  13'b0000110010011; // 403 0.09827443212270737
storage[5165] = -13'b0000000111010; // -58 -0.014148239977657795
storage[5166] = -13'b0000011111000; // -248 -0.06044871360063553
storage[5167] =  13'b0000001110001; // 113 0.027543693780899048
storage[5168] =  13'b0000010000110; // 134 0.03279704973101616
storage[5169] =  13'b0000001111011; // 123 0.03010687045753002
storage[5170] = -13'b0000110001111; // -399 -0.09738046675920486
storage[5171] =  13'b0000010111000; // 184 0.044986873865127563
storage[5172] =  13'b0000101110111; // 375 0.09159363806247711
storage[5173] =  13'b0000011000001; // 193 0.04708115756511688
storage[5174] =  13'b0000001001100; // 76 0.01864217035472393
storage[5175] =  13'b0000010001111; // 143 0.03480421006679535
storage[5176] = -13'b0000000001010; // -10 -0.0023532204795628786
storage[5177] =  13'b0000100111001; // 313 0.07640177756547928
storage[5178] = -13'b0011101011101; // -1885 -0.4600915312767029
storage[5179] =  13'b0001001100000; // 608 0.14847633242607117
storage[5180] =  13'b0000101000100; // 324 0.07904917001724243
storage[5181] =  13'b0000001110011; // 115 0.027984794229269028
storage[5182] =  13'b0000101100101; // 357 0.08704148977994919
storage[5183] = -13'b0000011010000; // -208 -0.05075477808713913
storage[5184] = -13'b0000011011110; // -222 -0.054158300161361694
storage[5185] =  13'b0000011000011; // 195 0.04751361161470413
storage[5186] =  13'b0000111011000; // 472 0.11520853638648987
storage[5187] = -13'b0000101110110; // -374 -0.09124589711427689
storage[5188] =  13'b0000100000000; // 256 0.0625174269080162
storage[5189] =  13'b0000010101110; // 174 0.042553313076496124
storage[5190] = -13'b0000010010100; // -148 -0.03603624179959297
storage[5191] =  13'b0000001011101; // 93 0.02259129285812378
storage[5192] =  13'b0000010011010; // 154 0.037687502801418304
storage[5193] =  13'b0000000100110; // 38 0.00921937171369791
storage[5194] =  13'b0000001011110; // 94 0.023064587265253067
storage[5195] =  13'b0000110110011; // 435 0.10629158467054367
storage[5196] =  13'b0000001000000; // 64 0.015739673748612404
storage[5197] =  13'b0000010010110; // 150 0.036692969501018524
storage[5198] = -13'b0000001000111; // -71 -0.017359759658575058
storage[5199] = -13'b0000010011111; // -159 -0.03884837403893471
storage[5200] =  13'b0000100011100; // 284 0.0693153515458107
storage[5201] = -13'b0000000001101; // -13 -0.0030569816008210182
storage[5202] =  13'b0000001000011; // 67 0.016351979225873947
storage[5203] = -13'b0000011100100; // -228 -0.055678777396678925
storage[5204] =  13'b0000011100100; // 228 0.05571594461798668
storage[5205] =  13'b0000100101001; // 297 0.07241054624319077
storage[5206] = -13'b0000000011001; // -25 -0.005985108204185963
storage[5207] =  13'b0000001110000; // 112 0.0273827463388443
storage[5208] =  13'b0000010111101; // 189 0.04606832563877106
storage[5209] =  13'b0000011100110; // 230 0.05616084486246109
storage[5210] =  13'b0000010110011; // 179 0.04378489404916763
storage[5211] = -13'b0000010001010; // -138 -0.03370102494955063
storage[5212] = -13'b0000001010000; // -80 -0.019418401643633842
storage[5213] =  13'b0000000010001; // 17 0.00427053589373827
storage[5214] = -13'b0000001101100; // -108 -0.026356030255556107
storage[5215] =  13'b0000100000100; // 260 0.0635647252202034
storage[5216] = -13'b0000001101110; // -110 -0.026806961745023727
storage[5217] = -13'b0000111100010; // -482 -0.11766031384468079
storage[5218] = -13'b0000000000111; // -7 -0.001755581353791058
storage[5219] = -13'b0000011100111; // -231 -0.05636833235621452
storage[5220] =  13'b0000001100101; // 101 0.024650106206536293
storage[5221] = -13'b0000000010011; // -19 -0.00475646834820509
storage[5222] =  13'b0000001110010; // 114 0.027789903804659843
storage[5223] =  13'b0000000011110; // 30 0.0072899856604635715
storage[5224] =  13'b0000011000010; // 194 0.04731030389666557
storage[5225] =  13'b0000100001110; // 270 0.0658869594335556
storage[5226] =  13'b0000000001011; // 11 0.002781103365123272
storage[5227] =  13'b0000100100001; // 289 0.0705464705824852
storage[5228] =  13'b0000010100110; // 166 0.04061891883611679
storage[5229] = -13'b0000000110100; // -52 -0.012791918590664864
storage[5230] = -13'b0000101110110; // -374 -0.09142125397920609
storage[5231] = -13'b0000111101110; // -494 -0.12055890262126923
storage[5232] = -13'b0000111000011; // -451 -0.11010672897100449
storage[5233] = -13'b0000010000101; // -133 -0.03238184005022049
storage[5234] =  13'b0000100001100; // 268 0.06537410616874695
storage[5235] =  13'b0000010111001; // 185 0.045128364115953445
storage[5236] = -13'b0000000110010; // -50 -0.012210221029818058
storage[5237] =  13'b0000100000001; // 257 0.06284681707620621
storage[5238] =  13'b0000000010001; // 17 0.004067813977599144
storage[5239] = -13'b0000111000010; // -450 -0.10987677425146103
storage[5240] = -13'b0000000110001; // -49 -0.012052168138325214
storage[5241] =  13'b0000011001011; // 203 0.049481648951768875
storage[5242] = -13'b0000000110011; // -51 -0.012469861656427383
storage[5243] =  13'b0000011010110; // 214 0.052173689007759094
storage[5244] = -13'b0000010010101; // -149 -0.0363512821495533
storage[5245] =  13'b0000001111100; // 124 0.030249010771512985
storage[5246] = -13'b0000000100110; // -38 -0.009344656951725483
storage[5247] =  13'b0000010001000; // 136 0.03319258242845535
storage[5248] = -13'b0000111011101; // -477 -0.1163514032959938
storage[5249] =  13'b0000000101010; // 42 0.010226646438241005
storage[5250] = -13'b0000100101011; // -299 -0.07305815070867538
storage[5251] = -13'b0001011011010; // -730 -0.17826221883296967
storage[5252] =  13'b0000110011100; // 412 0.10054566711187363
storage[5253] =  13'b0000001001111; // 79 0.019186383113265038
storage[5254] =  13'b0000110110111; // 439 0.10720814764499664
storage[5255] =  13'b0000100011000; // 280 0.06828789412975311
storage[5256] = -13'b0000110001010; // -394 -0.09626422822475433
storage[5257] = -13'b0000110011111; // -415 -0.10121691226959229
storage[5258] = -13'b0000000001000; // -8 -0.0018842363497242332
storage[5259] =  13'b0000011000010; // 194 0.04725100100040436
storage[5260] = -13'b0000001001010; // -74 -0.01811462827026844
storage[5261] =  13'b0000000111011; // 59 0.014451743103563786
storage[5262] =  13'b0000000000011; // 3 0.0006927614449523389
storage[5263] =  13'b0000001001001; // 73 0.01775301620364189
storage[5264] = -13'b0000001011110; // -94 -0.02301621250808239
storage[5265] =  13'b0000001011100; // 92 0.022454429417848587
storage[5266] = -13'b0001011110010; // -754 -0.18399780988693237
storage[5267] = -13'b0001000011001; // -537 -0.13108260929584503
storage[5268] = -13'b0000010010000; // -144 -0.03512407839298248
storage[5269] =  13'b0000000100100; // 36 0.008691789582371712
storage[5270] = -13'b0000101000010; // -322 -0.07865588366985321
storage[5271] = -13'b0000010001001; // -137 -0.033490151166915894
storage[5272] =  13'b0000000110000; // 48 0.011675504967570305
storage[5273] =  13'b0000010101000; // 168 0.04093789681792259
storage[5274] =  13'b0000100011001; // 281 0.06856530159711838
storage[5275] = -13'b0000110011001; // -409 -0.09974288195371628
storage[5276] = -13'b0000111111100; // -508 -0.12397277355194092
storage[5277] = -13'b0000001100101; // -101 -0.024567652493715286
storage[5278] = -13'b0000011110101; // -245 -0.05988585576415062
storage[5279] = -13'b0001011111001; // -761 -0.18576522171497345
storage[5280] =  13'b0000001000001; // 65 0.015761911869049072
storage[5281] =  13'b0000000101100; // 44 0.010845264419913292
storage[5282] = -13'b0000010100101; // -165 -0.040350452065467834
storage[5283] =  13'b0000000111011; // 59 0.01450777892023325
storage[5284] = -13'b0001000011111; // -543 -0.13262532651424408
storage[5285] =  13'b0001001110010; // 626 0.15284761786460876
storage[5286] = -13'b0001010000011; // -643 -0.15708401799201965
storage[5287] = -13'b0000110110110; // -438 -0.10698681324720383
storage[5288] = -13'b0000000101011; // -43 -0.01049697957932949
storage[5289] = -13'b0001011100011; // -739 -0.18039435148239136
storage[5290] = -13'b0000000011110; // -30 -0.007434620056301355
storage[5291] =  13'b0000001110100; // 116 0.028328128159046173
storage[5292] = -13'b0001101100000; // -864 -0.21097439527511597
storage[5293] =  13'b0001101101101; // 877 0.2141871154308319
storage[5294] =  13'b0000001111000; // 120 0.029334064573049545
storage[5295] =  13'b0001010101111; // 687 0.16775281727313995
storage[5296] =  13'b0001000000010; // 514 0.1254235804080963
storage[5297] = -13'b0001100110011; // -819 -0.1998872309923172
storage[5298] =  13'b0001010001001; // 649 0.15842947363853455
storage[5299] =  13'b0001001010111; // 599 0.14615003764629364
storage[5300] = -13'b0001011101101; // -749 -0.18291647732257843
storage[5301] = -13'b0001101011011; // -859 -0.20979149639606476
storage[5302] =  13'b0000110011000; // 408 0.09956136345863342
storage[5303] = -13'b0001010111000; // -696 -0.16997024416923523
storage[5304] = -13'b0001010100010; // -674 -0.16449590027332306
storage[5305] =  13'b0000000100000; // 32 0.007735949940979481
storage[5306] =  13'b0010000100000; // 1056 0.25776395201683044
storage[5307] =  13'b0000111101000; // 488 0.11915572732686996
storage[5308] =  13'b0000000010011; // 19 0.0047331303358078
storage[5309] = -13'b0001011010011; // -723 -0.1764049381017685
storage[5310] =  13'b0000111000111; // 455 0.11102302372455597
storage[5311] = -13'b0001011010010; // -722 -0.1763862818479538
storage[5312] =  13'b0010000110000; // 1072 0.26172396540641785
storage[5313] = -13'b0001010011010; // -666 -0.16256658732891083
storage[5314] = -13'b0001001110111; // -631 -0.1539759635925293
storage[5315] =  13'b0000011000011; // 195 0.04759177938103676
storage[5316] =  13'b0000011111001; // 249 0.06082851067185402
storage[5317] =  13'b0001011010001; // 721 0.1759837418794632
storage[5318] =  13'b0001100101100; // 812 0.19832992553710938
storage[5319] = -13'b0000111011111; // -479 -0.11688172072172165
storage[5320] = -13'b0000001111110; // -126 -0.030875451862812042
storage[5321] = -13'b0000010101110; // -174 -0.04253686964511871
storage[5322] = -13'b0000001100111; // -103 -0.025162428617477417
storage[5323] =  13'b0000100010110; // 278 0.06797172874212265
storage[5324] = -13'b0000100010010; // -274 -0.06681384146213531
storage[5325] = -13'b0000101100111; // -359 -0.08755665272474289
storage[5326] =  13'b0010100001101; // 1293 0.3156096637248993
storage[5327] = -13'b0000010000010; // -130 -0.03161768242716789
storage[5328] = -13'b0001011110100; // -756 -0.18444861471652985
storage[5329] =  13'b0000001001111; // 79 0.019265353679656982
storage[5330] = -13'b0001110111111; // -959 -0.23423956334590912
storage[5331] =  13'b0000010000010; // 130 0.03163379058241844
storage[5332] =  13'b0010101101011; // 1387 0.338686466217041
storage[5333] =  13'b0000000010001; // 17 0.0041803959757089615
storage[5334] =  13'b0000000010011; // 19 0.004748250357806683
storage[5335] = -13'b0000100111100; // -316 -0.07713864743709564
storage[5336] = -13'b0000000111011; // -59 -0.014432914555072784
storage[5337] =  13'b0000100100101; // 293 0.07149328291416168
storage[5338] =  13'b0001111010110; // 982 0.2398625910282135
storage[5339] = -13'b0000111110111; // -503 -0.1229059174656868
storage[5340] = -13'b0000101101100; // -364 -0.08875849097967148
storage[5341] = -13'b0001001001110; // -590 -0.14413423836231232
storage[5342] =  13'b0000001111101; // 125 0.030587663874030113
storage[5343] =  13'b0001100110001; // 817 0.199546217918396
storage[5344] = -13'b0000011111111; // -255 -0.06214180961251259
storage[5345] =  13'b0000001001110; // 78 0.018991755321621895
storage[5346] = -13'b0000001100010; // -98 -0.023857546970248222
storage[5347] = -13'b0000110001111; // -399 -0.09752011299133301
storage[5348] = -13'b0001000000111; // -519 -0.12661266326904297
storage[5349] = -13'b0000001000100; // -68 -0.016553835943341255
storage[5350] = -13'b0000100100101; // -293 -0.07147807627916336
storage[5351] =  13'b0010010110010; // 1202 0.2935124635696411
storage[5352] = -13'b0001010101100; // -684 -0.16697868704795837
storage[5353] = -13'b0000100101011; // -299 -0.07303519546985626
storage[5354] = -13'b0000100100010; // -290 -0.07077687978744507
storage[5355] =  13'b0000011110001; // 241 0.05879601463675499
storage[5356] =  13'b0000110011001; // 409 0.09978219866752625
storage[5357] =  13'b0001000100100; // 548 0.13386203348636627
storage[5358] = -13'b0000001001111; // -79 -0.019309554249048233
storage[5359] = -13'b0001111101010; // -1002 -0.24470099806785583
storage[5360] =  13'b0001010011011; // 667 0.16278918087482452
storage[5361] =  13'b0001000101101; // 557 0.13590845465660095
storage[5362] = -13'b0000111111001; // -505 -0.1232893243432045
storage[5363] = -13'b0000110011010; // -410 -0.10001981258392334
storage[5364] =  13'b0000111111101; // 509 0.12416382133960724
storage[5365] = -13'b0000001110110; // -118 -0.02882489003241062
storage[5366] = -13'b0000100001001; // -265 -0.06462208926677704
storage[5367] = -13'b0000100100010; // -290 -0.07088366895914078
storage[5368] =  13'b0001101111000; // 888 0.21686922013759613
storage[5369] = -13'b0000001011010; // -90 -0.02191053330898285
storage[5370] = -13'b0000110101100; // -428 -0.10456176102161407
storage[5371] = -13'b0001000111110; // -574 -0.14013637602329254
storage[5372] =  13'b0000011101010; // 234 0.05703065171837807
storage[5373] = -13'b0000100010100; // -276 -0.06746095418930054
storage[5374] = -13'b0000001101010; // -106 -0.02597091533243656
storage[5375] =  13'b0001110011001; // 921 0.22488248348236084
storage[5376] =  13'b0001010001001; // 649 0.15844228863716125
storage[5377] =  13'b0001000000001; // 513 0.12533697485923767
storage[5378] = -13'b0000011011100; // -220 -0.053767185658216476
storage[5379] =  13'b0000110111001; // 441 0.10756146907806396
storage[5380] =  13'b0000111011111; // 479 0.1170092225074768
storage[5381] =  13'b0000110000011; // 387 0.09451122581958771
storage[5382] = -13'b0000000011000; // -24 -0.005935312248766422
storage[5383] = -13'b0001000011110; // -542 -0.13239599764347076
storage[5384] = -13'b0000010010111; // -151 -0.03681783005595207
storage[5385] = -13'b0001011001001; // -713 -0.1741630584001541
storage[5386] = -13'b0000011100101; // -229 -0.05600607022643089
storage[5387] = -13'b0000001100010; // -98 -0.023886991664767265
storage[5388] =  13'b0010001110011; // 1139 0.27818092703819275
storage[5389] =  13'b0010000000000; // 1024 0.24990685284137726
storage[5390] = -13'b0001000101001; // -553 -0.13490994274616241
storage[5391] =  13'b0001100100001; // 801 0.19559694826602936
storage[5392] =  13'b0000101000110; // 326 0.07964883744716644
storage[5393] = -13'b0001101010000; // -848 -0.20709089934825897
storage[5394] = -13'b0010101110001; // -1393 -0.340060830116272
storage[5395] =  13'b0001001100010; // 610 0.1490303874015808
storage[5396] = -13'b0001010111111; // -703 -0.17152734100818634
storage[5397] =  13'b0001000110110; // 566 0.13823753595352173
storage[5398] =  13'b0001000110010; // 562 0.1371232122182846
storage[5399] =  13'b0000011111010; // 250 0.061019379645586014
storage[5400] =  13'b0001100000100; // 772 0.18855464458465576
storage[5401] = -13'b0000111001001; // -457 -0.11147185415029526
storage[5402] =  13'b0001011101101; // 749 0.182969331741333
storage[5403] =  13'b0000010000101; // 133 0.03234972432255745
storage[5404] = -13'b0000101011010; // -346 -0.08445696532726288
storage[5405] = -13'b0001101000100; // -836 -0.2041446566581726
storage[5406] = -13'b0000100100111; // -295 -0.07196313887834549
storage[5407] = -13'b0010010010111; // -1175 -0.28680554032325745
storage[5408] =  13'b0000000111100; // 60 0.014562501572072506
storage[5409] =  13'b0000101110100; // 372 0.09070633351802826
storage[5410] =  13'b0000011011100; // 220 0.053618308156728745
storage[5411] = -13'b0001100100111; // -807 -0.19708319008350372
storage[5412] =  13'b0001101001110; // 846 0.20653952658176422
storage[5413] =  13'b0000111001001; // 457 0.1115732192993164
storage[5414] =  13'b0001100010000; // 784 0.1913800686597824
storage[5415] =  13'b0001110010000; // 912 0.22276002168655396
storage[5416] =  13'b0000000110101; // 53 0.012900689616799355
storage[5417] =  13'b0000101011101; // 349 0.0852758139371872
storage[5418] =  13'b0000000010100; // 20 0.004846353083848953
storage[5419] = -13'b0001000001100; // -524 -0.12793339788913727
storage[5420] = -13'b0000111010111; // -471 -0.11508467048406601
storage[5421] = -13'b0000101110001; // -369 -0.090147003531456
storage[5422] = -13'b0001000110010; // -562 -0.13711799681186676
storage[5423] =  13'b0001010101100; // 684 0.16698971390724182
storage[5424] =  13'b0000100110001; // 305 0.07454967498779297
storage[5425] = -13'b0001100001110; // -782 -0.19084875285625458
storage[5426] = -13'b0010000000111; // -1031 -0.2518107295036316
storage[5427] =  13'b0000010010111; // 151 0.03690536320209503
storage[5428] = -13'b0000101111100; // -380 -0.09283263981342316
storage[5429] =  13'b0000110001001; // 393 0.09588854014873505
storage[5430] = -13'b0001100011110; // -798 -0.19487036764621735
storage[5431] =  13'b0001011000011; // 707 0.17253445088863373
storage[5432] =  13'b0000000000101; // 5 0.001177320722490549
storage[5433] =  13'b0000010001010; // 138 0.03371238335967064
storage[5434] =  13'b0001001000000; // 576 0.1407114565372467
storage[5435] = -13'b0001001111100; // -636 -0.15538464486598969
storage[5436] = -13'b0001000110101; // -565 -0.13790550827980042
storage[5437] =  13'b0000110101000; // 424 0.10358548909425735
storage[5438] = -13'b0001100000111; // -775 -0.1892244964838028
storage[5439] = -13'b0001011100110; // -742 -0.1811719536781311
storage[5440] = -13'b0000000111000; // -56 -0.013763817958533764
storage[5441] =  13'b0001010101010; // 682 0.1666223704814911
storage[5442] = -13'b0000000000110; // -6 -0.0015702510718256235
storage[5443] =  13'b0001100000110; // 774 0.18890225887298584
storage[5444] = -13'b0001101101110; // -878 -0.2142651230096817
storage[5445] = -13'b0110011111101; // -3325 -0.8117144703865051
storage[5446] = -13'b0001010111010; // -698 -0.17047716677188873
storage[5447] = -13'b0001101010010; // -850 -0.20752622187137604
storage[5448] =  13'b0000100001001; // 265 0.06462334841489792
storage[5449] =  13'b0111010001100; // 3724 0.9090909361839294
storage[5450] = -13'b0010010010000; // -1168 -0.2852747142314911
storage[5451] =  13'b0010101010101; // 1365 0.33320581912994385
storage[5452] = -13'b0011100001101; // -1805 -0.4406297206878662
storage[5453] =  13'b0011111011101; // 2013 0.4914056062698364
storage[5454] =  13'b0001000101010; // 554 0.13531462848186493
storage[5455] = -13'b0001110100011; // -931 -0.22736206650733948
storage[5456] = -13'b0011110101100; // -1964 -0.4795781672000885
storage[5457] = -13'b0110001011010; // -3162 -0.7719171643257141
storage[5458] = -13'b0001100011011; // -795 -0.1940820962190628
storage[5459] = -13'b0100010100100; // -2212 -0.5401360392570496



end

always @(posedge clk) if (we==1) storage[address_p] <= dp;
always @(posedge clk) if (re==1) datata<=storage[address];

endmodule
