module test();

parameter SIZE=12;

  reg clk;
  reg GO;
  reg signed [SIZE-1:0] storage [0:783]; 
  
  reg we_database;
  reg [SIZE-1:0] dp_database;
  reg [12:0] address_p_database;
  
  reg [9:0] x;
  
  wire [3:0] RESULT;
  TOP TOP(
	.clk					(clk),
	.GO						(GO),
	.RESULT					(RESULT),
	.we_database			(we_database), 
	.dp_database			(dp_database), 
	.address_p_database		(address_p_database-1), 
	.STOP					(STOP)
  );
initial begin
  clk=0;
  address_p_database=0;
  x=0;
  we_database=1;
  #200 GO=1;
end
always #10 clk=~clk;
always @(posedge clk)
	begin
		if (we_database)
		begin
			if (address_p_database<=783) 
				begin
						dp_database = storage[address_p_database];
						address_p_database=address_p_database+1'b1;
				end
			else we_database=0;
		end
		if ((x<=28*28)&&(GO)) x=x+1;
		else GO=0;
	if (STOP==1)
	begin
		$display("RESULT: %d",RESULT);
		$finish;
	end
 end
 
initial
	begin
		storage[0] =  11'b10011110000; // [0.6171875]
		storage[1] =  11'b10011111000; // [0.62109375]
		storage[2] =  11'b10100000000; // [0.625]
		storage[3] =  11'b10100010000; // [0.6328125]
		storage[4] =  11'b10100011000; // [0.63671875]
		storage[5] =  11'b10100011000; // [0.63671875]
		storage[6] =  11'b10100001000; // [0.62890625]
		storage[7] =  11'b10011010000; // [0.6015625]
		storage[8] =  11'b10001011000; // [0.54296875]
		storage[9] =  11'b01111011000; // [0.48046875]
		storage[10] =  11'b01101011000; // [0.41796875]
		storage[11] =  11'b01100100000; // [0.390625]
		storage[12] =  11'b01100011000; // [0.38671875]
		storage[13] =  11'b01101000000; // [0.40625]
		storage[14] =  11'b01110000000; // [0.4375]
		storage[15] =  11'b10000001000; // [0.50390625]
		storage[16] =  11'b10010101000; // [0.58203125]
		storage[17] =  11'b10100001000; // [0.62890625]
		storage[18] =  11'b10100101000; // [0.64453125]
		storage[19] =  11'b10100101000; // [0.64453125]
		storage[20] =  11'b10100110000; // [0.6484375]
		storage[21] =  11'b10100100000; // [0.640625]
		storage[22] =  11'b10100100000; // [0.640625]
		storage[23] =  11'b10100011000; // [0.63671875]
		storage[24] =  11'b10100010000; // [0.6328125]
		storage[25] =  11'b10100001000; // [0.62890625]
		storage[26] =  11'b10100000000; // [0.625]
		storage[27] =  11'b10011110000; // [0.6171875]
		storage[28] =  11'b10011101000; // [0.61328125]
		storage[29] =  11'b10011111000; // [0.62109375]
		storage[30] =  11'b10100000000; // [0.625]
		storage[31] =  11'b10100010000; // [0.6328125]
		storage[32] =  11'b10100011000; // [0.63671875]
		storage[33] =  11'b10100001000; // [0.62890625]
		storage[34] =  11'b10010110000; // [0.5859375]
		storage[35] =  11'b01110010000; // [0.4453125]
		storage[36] =  11'b01010010000; // [0.3203125]
		storage[37] =  11'b01000111000; // [0.27734375]
		storage[38] =  11'b01000011000; // [0.26171875]
		storage[39] =  11'b01000111000; // [0.27734375]
		storage[40] =  11'b01000111000; // [0.27734375]
		storage[41] =  11'b01000111000; // [0.27734375]
		storage[42] =  11'b01000111000; // [0.27734375]
		storage[43] =  11'b01010100000; // [0.328125]
		storage[44] =  11'b01110110000; // [0.4609375]
		storage[45] =  11'b10010111000; // [0.58984375]
		storage[46] =  11'b10100010000; // [0.6328125]
		storage[47] =  11'b10100101000; // [0.64453125]
		storage[48] =  11'b10100101000; // [0.64453125]
		storage[49] =  11'b10100100000; // [0.640625]
		storage[50] =  11'b10100101000; // [0.64453125]
		storage[51] =  11'b10100011000; // [0.63671875]
		storage[52] =  11'b10100011000; // [0.63671875]
		storage[53] =  11'b10100001000; // [0.62890625]
		storage[54] =  11'b10100000000; // [0.625]
		storage[55] =  11'b10011110000; // [0.6171875]
		storage[56] =  11'b10011100000; // [0.609375]
		storage[57] =  11'b10011110000; // [0.6171875]
		storage[58] =  11'b10100000000; // [0.625]
		storage[59] =  11'b10100001000; // [0.62890625]
		storage[60] =  11'b10100000000; // [0.625]
		storage[61] =  11'b10011001000; // [0.59765625]
		storage[62] =  11'b01110111000; // [0.46484375]
		storage[63] =  11'b01001010000; // [0.2890625]
		storage[64] =  11'b00111111000; // [0.24609375]
		storage[65] =  11'b01010000000; // [0.3125]
		storage[66] =  11'b01101101000; // [0.42578125]
		storage[67] =  11'b01111011000; // [0.48046875]
		storage[68] =  11'b01110001000; // [0.44140625]
		storage[69] =  11'b01011001000; // [0.34765625]
		storage[70] =  11'b01001000000; // [0.28125]
		storage[71] =  11'b01000011000; // [0.26171875]
		storage[72] =  11'b01010110000; // [0.3359375]
		storage[73] =  11'b01111111000; // [0.49609375]
		storage[74] =  11'b10011100000; // [0.609375]
		storage[75] =  11'b10100011000; // [0.63671875]
		storage[76] =  11'b10100100000; // [0.640625]
		storage[77] =  11'b10100101000; // [0.64453125]
		storage[78] =  11'b10100100000; // [0.640625]
		storage[79] =  11'b10100011000; // [0.63671875]
		storage[80] =  11'b10100010000; // [0.6328125]
		storage[81] =  11'b10100001000; // [0.62890625]
		storage[82] =  11'b10100000000; // [0.625]
		storage[83] =  11'b10011111000; // [0.62109375]
		storage[84] =  11'b10011101000; // [0.61328125]
		storage[85] =  11'b10011110000; // [0.6171875]
		storage[86] =  11'b10011111000; // [0.62109375]
		storage[87] =  11'b10011111000; // [0.62109375]
		storage[88] =  11'b10011011000; // [0.60546875]
		storage[89] =  11'b10000100000; // [0.515625]
		storage[90] =  11'b01001111000; // [0.30859375]
		storage[91] =  11'b00111111000; // [0.24609375]
		storage[92] =  11'b01010101000; // [0.33203125]
		storage[93] =  11'b10000001000; // [0.50390625]
		storage[94] =  11'b10011100000; // [0.609375]
		storage[95] =  11'b10100001000; // [0.62890625]
		storage[96] =  11'b10011100000; // [0.609375]
		storage[97] =  11'b10000111000; // [0.52734375]
		storage[98] =  11'b01100100000; // [0.390625]
		storage[99] =  11'b01001010000; // [0.2890625]
		storage[100] =  11'b01001001000; // [0.28515625]
		storage[101] =  11'b01101001000; // [0.41015625]
		storage[102] =  11'b10010000000; // [0.5625]
		storage[103] =  11'b10100000000; // [0.625]
		storage[104] =  11'b10100011000; // [0.63671875]
		storage[105] =  11'b10100101000; // [0.64453125]
		storage[106] =  11'b10100100000; // [0.640625]
		storage[107] =  11'b10100100000; // [0.640625]
		storage[108] =  11'b10100010000; // [0.6328125]
		storage[109] =  11'b10100001000; // [0.62890625]
		storage[110] =  11'b10100000000; // [0.625]
		storage[111] =  11'b10011111000; // [0.62109375]
		storage[112] =  11'b10011101000; // [0.61328125]
		storage[113] =  11'b10011101000; // [0.61328125]
		storage[114] =  11'b10011110000; // [0.6171875]
		storage[115] =  11'b10011101000; // [0.61328125]
		storage[116] =  11'b10010000000; // [0.5625]
		storage[117] =  11'b01011100000; // [0.359375]
		storage[118] =  11'b01000000000; // [0.25]
		storage[119] =  11'b01001011000; // [0.29296875]
		storage[120] =  11'b01111011000; // [0.48046875]
		storage[121] =  11'b10011110000; // [0.6171875]
		storage[122] =  11'b10100101000; // [0.64453125]
		storage[123] =  11'b10100111000; // [0.65234375]
		storage[124] =  11'b10101000000; // [0.65625]
		storage[125] =  11'b10011101000; // [0.61328125]
		storage[126] =  11'b10000001000; // [0.50390625]
		storage[127] =  11'b01011011000; // [0.35546875]
		storage[128] =  11'b01001010000; // [0.2890625]
		storage[129] =  11'b01010111000; // [0.33984375]
		storage[130] =  11'b10000010000; // [0.5078125]
		storage[131] =  11'b10011100000; // [0.609375]
		storage[132] =  11'b10100010000; // [0.6328125]
		storage[133] =  11'b10100100000; // [0.640625]
		storage[134] =  11'b10100101000; // [0.64453125]
		storage[135] =  11'b10100100000; // [0.640625]
		storage[136] =  11'b10100011000; // [0.63671875]
		storage[137] =  11'b10100010000; // [0.6328125]
		storage[138] =  11'b10100000000; // [0.625]
		storage[139] =  11'b10011111000; // [0.62109375]
		storage[140] =  11'b10011101000; // [0.61328125]
		storage[141] =  11'b10011110000; // [0.6171875]
		storage[142] =  11'b10011101000; // [0.61328125]
		storage[143] =  11'b10011000000; // [0.59375]
		storage[144] =  11'b01111001000; // [0.47265625]
		storage[145] =  11'b01000111000; // [0.27734375]
		storage[146] =  11'b01000110000; // [0.2734375]
		storage[147] =  11'b01101100000; // [0.421875]
		storage[148] =  11'b10010111000; // [0.58984375]
		storage[149] =  11'b10100011000; // [0.63671875]
		storage[150] =  11'b10101000000; // [0.65625]
		storage[151] =  11'b10101100000; // [0.671875]
		storage[152] =  11'b10101010000; // [0.6640625]
		storage[153] =  11'b10101000000; // [0.65625]
		storage[154] =  11'b10011001000; // [0.59765625]
		storage[155] =  11'b01111011000; // [0.48046875]
		storage[156] =  11'b01011001000; // [0.34765625]
		storage[157] =  11'b01010011000; // [0.32421875]
		storage[158] =  11'b01110101000; // [0.45703125]
		storage[159] =  11'b10011000000; // [0.59375]
		storage[160] =  11'b10100011000; // [0.63671875]
		storage[161] =  11'b10100110000; // [0.6484375]
		storage[162] =  11'b10100110000; // [0.6484375]
		storage[163] =  11'b10100110000; // [0.6484375]
		storage[164] =  11'b10100101000; // [0.64453125]
		storage[165] =  11'b10100011000; // [0.63671875]
		storage[166] =  11'b10100001000; // [0.62890625]
		storage[167] =  11'b10011111000; // [0.62109375]
		storage[168] =  11'b10011101000; // [0.61328125]
		storage[169] =  11'b10011101000; // [0.61328125]
		storage[170] =  11'b10011100000; // [0.609375]
		storage[171] =  11'b10001111000; // [0.55859375]
		storage[172] =  11'b01011110000; // [0.3671875]
		storage[173] =  11'b01001000000; // [0.28125]
		storage[174] =  11'b01100010000; // [0.3828125]
		storage[175] =  11'b10010000000; // [0.5625]
		storage[176] =  11'b10100010000; // [0.6328125]
		storage[177] =  11'b10100111000; // [0.65234375]
		storage[178] =  11'b10101100000; // [0.671875]
		storage[179] =  11'b10101101000; // [0.67578125]
		storage[180] =  11'b10101100000; // [0.671875]
		storage[181] =  11'b10101011000; // [0.66796875]
		storage[182] =  11'b10100111000; // [0.65234375]
		storage[183] =  11'b10010100000; // [0.578125]
		storage[184] =  11'b01110001000; // [0.44140625]
		storage[185] =  11'b01010111000; // [0.33984375]
		storage[186] =  11'b01101101000; // [0.42578125]
		storage[187] =  11'b10010011000; // [0.57421875]
		storage[188] =  11'b10100010000; // [0.6328125]
		storage[189] =  11'b10101000000; // [0.65625]
		storage[190] =  11'b10101000000; // [0.65625]
		storage[191] =  11'b10101000000; // [0.65625]
		storage[192] =  11'b10100110000; // [0.6484375]
		storage[193] =  11'b10100100000; // [0.640625]
		storage[194] =  11'b10100010000; // [0.6328125]
		storage[195] =  11'b10011111000; // [0.62109375]
		storage[196] =  11'b10011101000; // [0.61328125]
		storage[197] =  11'b10011110000; // [0.6171875]
		storage[198] =  11'b10011001000; // [0.59765625]
		storage[199] =  11'b01111111000; // [0.49609375]
		storage[200] =  11'b01001110000; // [0.3046875]
		storage[201] =  11'b01010000000; // [0.3125]
		storage[202] =  11'b01111011000; // [0.48046875]
		storage[203] =  11'b10011111000; // [0.62109375]
		storage[204] =  11'b10100110000; // [0.6484375]
		storage[205] =  11'b10101011000; // [0.66796875]
		storage[206] =  11'b10101111000; // [0.68359375]
		storage[207] =  11'b10101111000; // [0.68359375]
		storage[208] =  11'b10101110000; // [0.6796875]
		storage[209] =  11'b10101101000; // [0.67578125]
		storage[210] =  11'b10101011000; // [0.66796875]
		storage[211] =  11'b10100000000; // [0.625]
		storage[212] =  11'b10000000000; // [0.5]
		storage[213] =  11'b01011101000; // [0.36328125]
		storage[214] =  11'b01101010000; // [0.4140625]
		storage[215] =  11'b10010000000; // [0.5625]
		storage[216] =  11'b10100010000; // [0.6328125]
		storage[217] =  11'b10101000000; // [0.65625]
		storage[218] =  11'b10101010000; // [0.6640625]
		storage[219] =  11'b10101000000; // [0.65625]
		storage[220] =  11'b10101000000; // [0.65625]
		storage[221] =  11'b10100100000; // [0.640625]
		storage[222] =  11'b10100011000; // [0.63671875]
		storage[223] =  11'b10100000000; // [0.625]
		storage[224] =  11'b10011110000; // [0.6171875]
		storage[225] =  11'b10011101000; // [0.61328125]
		storage[226] =  11'b10010101000; // [0.58203125]
		storage[227] =  11'b01101101000; // [0.42578125]
		storage[228] =  11'b01001000000; // [0.28125]
		storage[229] =  11'b01011101000; // [0.36328125]
		storage[230] =  11'b10001101000; // [0.55078125]
		storage[231] =  11'b10100011000; // [0.63671875]
		storage[232] =  11'b10101011000; // [0.66796875]
		storage[233] =  11'b10101110000; // [0.6796875]
		storage[234] =  11'b10110000000; // [0.6875]
		storage[235] =  11'b10110000000; // [0.6875]
		storage[236] =  11'b10110000000; // [0.6875]
		storage[237] =  11'b10101111000; // [0.68359375]
		storage[238] =  11'b10101100000; // [0.671875]
		storage[239] =  11'b10100101000; // [0.64453125]
		storage[240] =  11'b10001000000; // [0.53125]
		storage[241] =  11'b01100010000; // [0.3828125]
		storage[242] =  11'b01100101000; // [0.39453125]
		storage[243] =  11'b10001100000; // [0.546875]
		storage[244] =  11'b10100001000; // [0.62890625]
		storage[245] =  11'b10101001000; // [0.66015625]
		storage[246] =  11'b10101010000; // [0.6640625]
		storage[247] =  11'b10101011000; // [0.66796875]
		storage[248] =  11'b10100111000; // [0.65234375]
		storage[249] =  11'b10100110000; // [0.6484375]
		storage[250] =  11'b10100011000; // [0.63671875]
		storage[251] =  11'b10100000000; // [0.625]
		storage[252] =  11'b10011100000; // [0.609375]
		storage[253] =  11'b10011100000; // [0.609375]
		storage[254] =  11'b10001111000; // [0.55859375]
		storage[255] =  11'b01011111000; // [0.37109375]
		storage[256] =  11'b01001000000; // [0.28125]
		storage[257] =  11'b01101101000; // [0.42578125]
		storage[258] =  11'b10011011000; // [0.60546875]
		storage[259] =  11'b10100111000; // [0.65234375]
		storage[260] =  11'b10101101000; // [0.67578125]
		storage[261] =  11'b10110000000; // [0.6875]
		storage[262] =  11'b10110000000; // [0.6875]
		storage[263] =  11'b10110000000; // [0.6875]
		storage[264] =  11'b10110000000; // [0.6875]
		storage[265] =  11'b10110000000; // [0.6875]
		storage[266] =  11'b10101110000; // [0.6796875]
		storage[267] =  11'b10101000000; // [0.65625]
		storage[268] =  11'b10001100000; // [0.546875]
		storage[269] =  11'b01100110000; // [0.3984375]
		storage[270] =  11'b01011100000; // [0.359375]
		storage[271] =  11'b10000110000; // [0.5234375]
		storage[272] =  11'b10011111000; // [0.62109375]
		storage[273] =  11'b10101000000; // [0.65625]
		storage[274] =  11'b10101010000; // [0.6640625]
		storage[275] =  11'b10101001000; // [0.66015625]
		storage[276] =  11'b10101000000; // [0.65625]
		storage[277] =  11'b10100110000; // [0.6484375]
		storage[278] =  11'b10100010000; // [0.6328125]
		storage[279] =  11'b10100001000; // [0.62890625]
		storage[280] =  11'b10011100000; // [0.609375]
		storage[281] =  11'b10011010000; // [0.6015625]
		storage[282] =  11'b10000110000; // [0.5234375]
		storage[283] =  11'b01010011000; // [0.32421875]
		storage[284] =  11'b01001101000; // [0.30078125]
		storage[285] =  11'b01111010000; // [0.4765625]
		storage[286] =  11'b10100000000; // [0.625]
		storage[287] =  11'b10101000000; // [0.65625]
		storage[288] =  11'b10101110000; // [0.6796875]
		storage[289] =  11'b10101111000; // [0.68359375]
		storage[290] =  11'b10110000000; // [0.6875]
		storage[291] =  11'b10110000000; // [0.6875]
		storage[292] =  11'b10110001000; // [0.69140625]
		storage[293] =  11'b10110000000; // [0.6875]
		storage[294] =  11'b10101110000; // [0.6796875]
		storage[295] =  11'b10101001000; // [0.66015625]
		storage[296] =  11'b10001111000; // [0.55859375]
		storage[297] =  11'b01101000000; // [0.40625]
		storage[298] =  11'b01010111000; // [0.33984375]
		storage[299] =  11'b10000010000; // [0.5078125]
		storage[300] =  11'b10011110000; // [0.6171875]
		storage[301] =  11'b10100111000; // [0.65234375]
		storage[302] =  11'b10101010000; // [0.6640625]
		storage[303] =  11'b10101001000; // [0.66015625]
		storage[304] =  11'b10100111000; // [0.65234375]
		storage[305] =  11'b10100110000; // [0.6484375]
		storage[306] =  11'b10100010000; // [0.6328125]
		storage[307] =  11'b10100000000; // [0.625]
		storage[308] =  11'b10011101000; // [0.61328125]
		storage[309] =  11'b10011000000; // [0.59375]
		storage[310] =  11'b01111100000; // [0.484375]
		storage[311] =  11'b01001100000; // [0.296875]
		storage[312] =  11'b01010011000; // [0.32421875]
		storage[313] =  11'b10001001000; // [0.53515625]
		storage[314] =  11'b10100010000; // [0.6328125]
		storage[315] =  11'b10101010000; // [0.6640625]
		storage[316] =  11'b10101101000; // [0.67578125]
		storage[317] =  11'b10101110000; // [0.6796875]
		storage[318] =  11'b10101110000; // [0.6796875]
		storage[319] =  11'b10110000000; // [0.6875]
		storage[320] =  11'b10110000000; // [0.6875]
		storage[321] =  11'b10110000000; // [0.6875]
		storage[322] =  11'b10101110000; // [0.6796875]
		storage[323] =  11'b10101001000; // [0.66015625]
		storage[324] =  11'b10001110000; // [0.5546875]
		storage[325] =  11'b01101000000; // [0.40625]
		storage[326] =  11'b01010110000; // [0.3359375]
		storage[327] =  11'b10000000000; // [0.5]
		storage[328] =  11'b10011101000; // [0.61328125]
		storage[329] =  11'b10100110000; // [0.6484375]
		storage[330] =  11'b10101000000; // [0.65625]
		storage[331] =  11'b10101000000; // [0.65625]
		storage[332] =  11'b10100111000; // [0.65234375]
		storage[333] =  11'b10100100000; // [0.640625]
		storage[334] =  11'b10100001000; // [0.62890625]
		storage[335] =  11'b10011111000; // [0.62109375]
		storage[336] =  11'b10011100000; // [0.609375]
		storage[337] =  11'b10010100000; // [0.578125]
		storage[338] =  11'b01101111000; // [0.43359375]
		storage[339] =  11'b01000111000; // [0.27734375]
		storage[340] =  11'b01011100000; // [0.359375]
		storage[341] =  11'b10001111000; // [0.55859375]
		storage[342] =  11'b10100100000; // [0.640625]
		storage[343] =  11'b10101001000; // [0.66015625]
		storage[344] =  11'b10101100000; // [0.671875]
		storage[345] =  11'b10101100000; // [0.671875]
		storage[346] =  11'b10101101000; // [0.67578125]
		storage[347] =  11'b10101110000; // [0.6796875]
		storage[348] =  11'b10101110000; // [0.6796875]
		storage[349] =  11'b10101110000; // [0.6796875]
		storage[350] =  11'b10101011000; // [0.66796875]
		storage[351] =  11'b10100110000; // [0.6484375]
		storage[352] =  11'b10001101000; // [0.55078125]
		storage[353] =  11'b01100110000; // [0.3984375]
		storage[354] =  11'b01010101000; // [0.33203125]
		storage[355] =  11'b10000010000; // [0.5078125]
		storage[356] =  11'b10011101000; // [0.61328125]
		storage[357] =  11'b10100100000; // [0.640625]
		storage[358] =  11'b10101000000; // [0.65625]
		storage[359] =  11'b10100111000; // [0.65234375]
		storage[360] =  11'b10100101000; // [0.64453125]
		storage[361] =  11'b10100011000; // [0.63671875]
		storage[362] =  11'b10100001000; // [0.62890625]
		storage[363] =  11'b10011110000; // [0.6171875]
		storage[364] =  11'b10011010000; // [0.6015625]
		storage[365] =  11'b10010000000; // [0.5625]
		storage[366] =  11'b01100100000; // [0.390625]
		storage[367] =  11'b01000111000; // [0.27734375]
		storage[368] =  11'b01100110000; // [0.3984375]
		storage[369] =  11'b10010101000; // [0.58203125]
		storage[370] =  11'b10100011000; // [0.63671875]
		storage[371] =  11'b10101000000; // [0.65625]
		storage[372] =  11'b10101011000; // [0.66796875]
		storage[373] =  11'b10101011000; // [0.66796875]
		storage[374] =  11'b10101011000; // [0.66796875]
		storage[375] =  11'b10101100000; // [0.671875]
		storage[376] =  11'b10101101000; // [0.67578125]
		storage[377] =  11'b10101011000; // [0.66796875]
		storage[378] =  11'b10101001000; // [0.66015625]
		storage[379] =  11'b10100011000; // [0.63671875]
		storage[380] =  11'b10001010000; // [0.5390625]
		storage[381] =  11'b01100010000; // [0.3828125]
		storage[382] =  11'b01010111000; // [0.33984375]
		storage[383] =  11'b10000110000; // [0.5234375]
		storage[384] =  11'b10011110000; // [0.6171875]
		storage[385] =  11'b10100101000; // [0.64453125]
		storage[386] =  11'b10100101000; // [0.64453125]
		storage[387] =  11'b10100101000; // [0.64453125]
		storage[388] =  11'b10100100000; // [0.640625]
		storage[389] =  11'b10100010000; // [0.6328125]
		storage[390] =  11'b10100000000; // [0.625]
		storage[391] =  11'b10011110000; // [0.6171875]
		storage[392] =  11'b10011001000; // [0.59765625]
		storage[393] =  11'b10001100000; // [0.546875]
		storage[394] =  11'b01011111000; // [0.37109375]
		storage[395] =  11'b01000111000; // [0.27734375]
		storage[396] =  11'b01101100000; // [0.421875]
		storage[397] =  11'b10011000000; // [0.59375]
		storage[398] =  11'b10100100000; // [0.640625]
		storage[399] =  11'b10100111000; // [0.65234375]
		storage[400] =  11'b10101001000; // [0.66015625]
		storage[401] =  11'b10101010000; // [0.6640625]
		storage[402] =  11'b10101100000; // [0.671875]
		storage[403] =  11'b10101100000; // [0.671875]
		storage[404] =  11'b10101100000; // [0.671875]
		storage[405] =  11'b10101011000; // [0.66796875]
		storage[406] =  11'b10101001000; // [0.66015625]
		storage[407] =  11'b10011111000; // [0.62109375]
		storage[408] =  11'b10000000000; // [0.5]
		storage[409] =  11'b01010111000; // [0.33984375]
		storage[410] =  11'b01011010000; // [0.3515625]
		storage[411] =  11'b10001010000; // [0.5390625]
		storage[412] =  11'b10011111000; // [0.62109375]
		storage[413] =  11'b10100101000; // [0.64453125]
		storage[414] =  11'b10100101000; // [0.64453125]
		storage[415] =  11'b10100101000; // [0.64453125]
		storage[416] =  11'b10100011000; // [0.63671875]
		storage[417] =  11'b10100001000; // [0.62890625]
		storage[418] =  11'b10011111000; // [0.62109375]
		storage[419] =  11'b10011101000; // [0.61328125]
		storage[420] =  11'b10011001000; // [0.59765625]
		storage[421] =  11'b10001010000; // [0.5390625]
		storage[422] =  11'b01011111000; // [0.37109375]
		storage[423] =  11'b01001010000; // [0.2890625]
		storage[424] =  11'b01101101000; // [0.42578125]
		storage[425] =  11'b10011001000; // [0.59765625]
		storage[426] =  11'b10100011000; // [0.63671875]
		storage[427] =  11'b10100111000; // [0.65234375]
		storage[428] =  11'b10101000000; // [0.65625]
		storage[429] =  11'b10101001000; // [0.66015625]
		storage[430] =  11'b10101010000; // [0.6640625]
		storage[431] =  11'b10101010000; // [0.6640625]
		storage[432] =  11'b10101011000; // [0.66796875]
		storage[433] =  11'b10101011000; // [0.66796875]
		storage[434] =  11'b10101001000; // [0.66015625]
		storage[435] =  11'b10011010000; // [0.6015625]
		storage[436] =  11'b01110100000; // [0.453125]
		storage[437] =  11'b01001100000; // [0.296875]
		storage[438] =  11'b01011100000; // [0.359375]
		storage[439] =  11'b10001101000; // [0.55078125]
		storage[440] =  11'b10100000000; // [0.625]
		storage[441] =  11'b10100100000; // [0.640625]
		storage[442] =  11'b10100100000; // [0.640625]
		storage[443] =  11'b10100100000; // [0.640625]
		storage[444] =  11'b10100010000; // [0.6328125]
		storage[445] =  11'b10100000000; // [0.625]
		storage[446] =  11'b10011110000; // [0.6171875]
		storage[447] =  11'b10011101000; // [0.61328125]
		storage[448] =  11'b10011000000; // [0.59375]
		storage[449] =  11'b10001100000; // [0.546875]
		storage[450] =  11'b01100100000; // [0.390625]
		storage[451] =  11'b01001010000; // [0.2890625]
		storage[452] =  11'b01101001000; // [0.41015625]
		storage[453] =  11'b10010100000; // [0.578125]
		storage[454] =  11'b10100010000; // [0.6328125]
		storage[455] =  11'b10100100000; // [0.640625]
		storage[456] =  11'b10100111000; // [0.65234375]
		storage[457] =  11'b10100110000; // [0.6484375]
		storage[458] =  11'b10100111000; // [0.65234375]
		storage[459] =  11'b10101010000; // [0.6640625]
		storage[460] =  11'b10101010000; // [0.6640625]
		storage[461] =  11'b10101010000; // [0.6640625]
		storage[462] =  11'b10100111000; // [0.65234375]
		storage[463] =  11'b10001111000; // [0.55859375]
		storage[464] =  11'b01100010000; // [0.3828125]
		storage[465] =  11'b01000110000; // [0.2734375]
		storage[466] =  11'b01100010000; // [0.3828125]
		storage[467] =  11'b10010000000; // [0.5625]
		storage[468] =  11'b10100000000; // [0.625]
		storage[469] =  11'b10100011000; // [0.63671875]
		storage[470] =  11'b10100011000; // [0.63671875]
		storage[471] =  11'b10100010000; // [0.6328125]
		storage[472] =  11'b10100000000; // [0.625]
		storage[473] =  11'b10011111000; // [0.62109375]
		storage[474] =  11'b10011110000; // [0.6171875]
		storage[475] =  11'b10011100000; // [0.609375]
		storage[476] =  11'b10011010000; // [0.6015625]
		storage[477] =  11'b10010001000; // [0.56640625]
		storage[478] =  11'b01110001000; // [0.44140625]
		storage[479] =  11'b01001100000; // [0.296875]
		storage[480] =  11'b01100110000; // [0.3984375]
		storage[481] =  11'b10010010000; // [0.5703125]
		storage[482] =  11'b10100000000; // [0.625]
		storage[483] =  11'b10100101000; // [0.64453125]
		storage[484] =  11'b10100101000; // [0.64453125]
		storage[485] =  11'b10100111000; // [0.65234375]
		storage[486] =  11'b10101000000; // [0.65625]
		storage[487] =  11'b10101010000; // [0.6640625]
		storage[488] =  11'b10101011000; // [0.66796875]
		storage[489] =  11'b10101001000; // [0.66015625]
		storage[490] =  11'b10011110000; // [0.6171875]
		storage[491] =  11'b01111001000; // [0.47265625]
		storage[492] =  11'b01001101000; // [0.30078125]
		storage[493] =  11'b01000100000; // [0.265625]
		storage[494] =  11'b01110010000; // [0.4453125]
		storage[495] =  11'b10011000000; // [0.59375]
		storage[496] =  11'b10100011000; // [0.63671875]
		storage[497] =  11'b10100100000; // [0.640625]
		storage[498] =  11'b10100101000; // [0.64453125]
		storage[499] =  11'b10100011000; // [0.63671875]
		storage[500] =  11'b10100001000; // [0.62890625]
		storage[501] =  11'b10011111000; // [0.62109375]
		storage[502] =  11'b10011110000; // [0.6171875]
		storage[503] =  11'b10011101000; // [0.61328125]
		storage[504] =  11'b10011011000; // [0.60546875]
		storage[505] =  11'b10010100000; // [0.578125]
		storage[506] =  11'b01111101000; // [0.48828125]
		storage[507] =  11'b01010010000; // [0.3203125]
		storage[508] =  11'b01100010000; // [0.3828125]
		storage[509] =  11'b10001110000; // [0.5546875]
		storage[510] =  11'b10011111000; // [0.62109375]
		storage[511] =  11'b10100011000; // [0.63671875]
		storage[512] =  11'b10100101000; // [0.64453125]
		storage[513] =  11'b10100110000; // [0.6484375]
		storage[514] =  11'b10101000000; // [0.65625]
		storage[515] =  11'b10101010000; // [0.6640625]
		storage[516] =  11'b10101010000; // [0.6640625]
		storage[517] =  11'b10101000000; // [0.65625]
		storage[518] =  11'b10001101000; // [0.55078125]
		storage[519] =  11'b01011111000; // [0.37109375]
		storage[520] =  11'b01000000000; // [0.25]
		storage[521] =  11'b01001000000; // [0.28125]
		storage[522] =  11'b10000011000; // [0.51171875]
		storage[523] =  11'b10011101000; // [0.61328125]
		storage[524] =  11'b10100100000; // [0.640625]
		storage[525] =  11'b10100110000; // [0.6484375]
		storage[526] =  11'b10100011000; // [0.63671875]
		storage[527] =  11'b10100011000; // [0.63671875]
		storage[528] =  11'b10100001000; // [0.62890625]
		storage[529] =  11'b10011111000; // [0.62109375]
		storage[530] =  11'b10011110000; // [0.6171875]
		storage[531] =  11'b10011100000; // [0.609375]
		storage[532] =  11'b10011001000; // [0.59765625]
		storage[533] =  11'b10010101000; // [0.58203125]
		storage[534] =  11'b10000110000; // [0.5234375]
		storage[535] =  11'b01011110000; // [0.3671875]
		storage[536] =  11'b01010111000; // [0.33984375]
		storage[537] =  11'b10000010000; // [0.5078125]
		storage[538] =  11'b10011100000; // [0.609375]
		storage[539] =  11'b10100001000; // [0.62890625]
		storage[540] =  11'b10100011000; // [0.63671875]
		storage[541] =  11'b10100101000; // [0.64453125]
		storage[542] =  11'b10100110000; // [0.6484375]
		storage[543] =  11'b10101001000; // [0.66015625]
		storage[544] =  11'b10101001000; // [0.66015625]
		storage[545] =  11'b10011111000; // [0.62109375]
		storage[546] =  11'b01111100000; // [0.484375]
		storage[547] =  11'b01001011000; // [0.29296875]
		storage[548] =  11'b00111010000; // [0.2265625]
		storage[549] =  11'b01010010000; // [0.3203125]
		storage[550] =  11'b10001011000; // [0.54296875]
		storage[551] =  11'b10011111000; // [0.62109375]
		storage[552] =  11'b10100101000; // [0.64453125]
		storage[553] =  11'b10100011000; // [0.63671875]
		storage[554] =  11'b10100010000; // [0.6328125]
		storage[555] =  11'b10100000000; // [0.625]
		storage[556] =  11'b10011110000; // [0.6171875]
		storage[557] =  11'b10011101000; // [0.61328125]
		storage[558] =  11'b10011100000; // [0.609375]
		storage[559] =  11'b10011011000; // [0.60546875]
		storage[560] =  11'b10010111000; // [0.58984375]
		storage[561] =  11'b10010110000; // [0.5859375]
		storage[562] =  11'b10001101000; // [0.55078125]
		storage[563] =  11'b01101111000; // [0.43359375]
		storage[564] =  11'b01010100000; // [0.328125]
		storage[565] =  11'b01110010000; // [0.4453125]
		storage[566] =  11'b10010111000; // [0.58984375]
		storage[567] =  11'b10011111000; // [0.62109375]
		storage[568] =  11'b10100010000; // [0.6328125]
		storage[569] =  11'b10100011000; // [0.63671875]
		storage[570] =  11'b10100111000; // [0.65234375]
		storage[571] =  11'b10100111000; // [0.65234375]
		storage[572] =  11'b10101000000; // [0.65625]
		storage[573] =  11'b10010111000; // [0.58984375]
		storage[574] =  11'b01101101000; // [0.42578125]
		storage[575] =  11'b01000010000; // [0.2578125]
		storage[576] =  11'b00111010000; // [0.2265625]
		storage[577] =  11'b01100001000; // [0.37890625]
		storage[578] =  11'b10010011000; // [0.57421875]
		storage[579] =  11'b10100001000; // [0.62890625]
		storage[580] =  11'b10100101000; // [0.64453125]
		storage[581] =  11'b10100010000; // [0.6328125]
		storage[582] =  11'b10100000000; // [0.625]
		storage[583] =  11'b10011111000; // [0.62109375]
		storage[584] =  11'b10011110000; // [0.6171875]
		storage[585] =  11'b10011100000; // [0.609375]
		storage[586] =  11'b10011010000; // [0.6015625]
		storage[587] =  11'b10011001000; // [0.59765625]
		storage[588] =  11'b10010111000; // [0.58984375]
		storage[589] =  11'b10010111000; // [0.58984375]
		storage[590] =  11'b10010011000; // [0.57421875]
		storage[591] =  11'b10000010000; // [0.5078125]
		storage[592] =  11'b01011100000; // [0.359375]
		storage[593] =  11'b01100011000; // [0.38671875]
		storage[594] =  11'b10001010000; // [0.5390625]
		storage[595] =  11'b10011101000; // [0.61328125]
		storage[596] =  11'b10100001000; // [0.62890625]
		storage[597] =  11'b10100011000; // [0.63671875]
		storage[598] =  11'b10100100000; // [0.640625]
		storage[599] =  11'b10100101000; // [0.64453125]
		storage[600] =  11'b10011111000; // [0.62109375]
		storage[601] =  11'b10000000000; // [0.5]
		storage[602] =  11'b01010010000; // [0.3203125]
		storage[603] =  11'b00111001000; // [0.22265625]
		storage[604] =  11'b01000000000; // [0.25]
		storage[605] =  11'b01110110000; // [0.4609375]
		storage[606] =  11'b10011010000; // [0.6015625]
		storage[607] =  11'b10100010000; // [0.6328125]
		storage[608] =  11'b10100011000; // [0.63671875]
		storage[609] =  11'b10100001000; // [0.62890625]
		storage[610] =  11'b10100000000; // [0.625]
		storage[611] =  11'b10011111000; // [0.62109375]
		storage[612] =  11'b10011101000; // [0.61328125]
		storage[613] =  11'b10011011000; // [0.60546875]
		storage[614] =  11'b10011001000; // [0.59765625]
		storage[615] =  11'b10010111000; // [0.58984375]
		storage[616] =  11'b10010110000; // [0.5859375]
		storage[617] =  11'b10010110000; // [0.5859375]
		storage[618] =  11'b10010110000; // [0.5859375]
		storage[619] =  11'b10001101000; // [0.55078125]
		storage[620] =  11'b01110011000; // [0.44921875]
		storage[621] =  11'b01010101000; // [0.33203125]
		storage[622] =  11'b01101110000; // [0.4296875]
		storage[623] =  11'b10010000000; // [0.5625]
		storage[624] =  11'b10011100000; // [0.609375]
		storage[625] =  11'b10100000000; // [0.625]
		storage[626] =  11'b10100000000; // [0.625]
		storage[627] =  11'b10011110000; // [0.6171875]
		storage[628] =  11'b10001000000; // [0.53125]
		storage[629] =  11'b01011001000; // [0.34765625]
		storage[630] =  11'b00111010000; // [0.2265625]
		storage[631] =  11'b00111010000; // [0.2265625]
		storage[632] =  11'b01010101000; // [0.33203125]
		storage[633] =  11'b10001000000; // [0.53125]
		storage[634] =  11'b10011100000; // [0.609375]
		storage[635] =  11'b10100000000; // [0.625]
		storage[636] =  11'b10100000000; // [0.625]
		storage[637] =  11'b10011111000; // [0.62109375]
		storage[638] =  11'b10011101000; // [0.61328125]
		storage[639] =  11'b10011100000; // [0.609375]
		storage[640] =  11'b10011010000; // [0.6015625]
		storage[641] =  11'b10010111000; // [0.58984375]
		storage[642] =  11'b10010110000; // [0.5859375]
		storage[643] =  11'b10010101000; // [0.58203125]
		storage[644] =  11'b10010100000; // [0.578125]
		storage[645] =  11'b10010100000; // [0.578125]
		storage[646] =  11'b10010110000; // [0.5859375]
		storage[647] =  11'b10010011000; // [0.57421875]
		storage[648] =  11'b10000100000; // [0.515625]
		storage[649] =  11'b01011100000; // [0.359375]
		storage[650] =  11'b01001100000; // [0.296875]
		storage[651] =  11'b01100000000; // [0.375]
		storage[652] =  11'b01111110000; // [0.4921875]
		storage[653] =  11'b10010001000; // [0.56640625]
		storage[654] =  11'b10010011000; // [0.57421875]
		storage[655] =  11'b10000100000; // [0.515625]
		storage[656] =  11'b01011111000; // [0.37109375]
		storage[657] =  11'b00111110000; // [0.2421875]
		storage[658] =  11'b00111001000; // [0.22265625]
		storage[659] =  11'b01001101000; // [0.30078125]
		storage[660] =  11'b01111010000; // [0.4765625]
		storage[661] =  11'b10011000000; // [0.59375]
		storage[662] =  11'b10011110000; // [0.6171875]
		storage[663] =  11'b10011110000; // [0.6171875]
		storage[664] =  11'b10011110000; // [0.6171875]
		storage[665] =  11'b10011101000; // [0.61328125]
		storage[666] =  11'b10011100000; // [0.609375]
		storage[667] =  11'b10011010000; // [0.6015625]
		storage[668] =  11'b10011000000; // [0.59375]
		storage[669] =  11'b10010111000; // [0.58984375]
		storage[670] =  11'b10010110000; // [0.5859375]
		storage[671] =  11'b10010011000; // [0.57421875]
		storage[672] =  11'b10010011000; // [0.57421875]
		storage[673] =  11'b10010101000; // [0.58203125]
		storage[674] =  11'b10010110000; // [0.5859375]
		storage[675] =  11'b10010110000; // [0.5859375]
		storage[676] =  11'b10001111000; // [0.55859375]
		storage[677] =  11'b01110111000; // [0.46484375]
		storage[678] =  11'b01001011000; // [0.29296875]
		storage[679] =  11'b00111101000; // [0.23828125]
		storage[680] =  11'b01001000000; // [0.28125]
		storage[681] =  11'b01010100000; // [0.328125]
		storage[682] =  11'b01010101000; // [0.33203125]
		storage[683] =  11'b01001000000; // [0.28125]
		storage[684] =  11'b00111100000; // [0.234375]
		storage[685] =  11'b00111101000; // [0.23828125]
		storage[686] =  11'b01010010000; // [0.3203125]
		storage[687] =  11'b01111010000; // [0.4765625]
		storage[688] =  11'b10010111000; // [0.58984375]
		storage[689] =  11'b10011101000; // [0.61328125]
		storage[690] =  11'b10011110000; // [0.6171875]
		storage[691] =  11'b10011100000; // [0.609375]
		storage[692] =  11'b10011101000; // [0.61328125]
		storage[693] =  11'b10011100000; // [0.609375]
		storage[694] =  11'b10011010000; // [0.6015625]
		storage[695] =  11'b10011001000; // [0.59765625]
		storage[696] =  11'b10010111000; // [0.58984375]
		storage[697] =  11'b10010110000; // [0.5859375]
		storage[698] =  11'b10010101000; // [0.58203125]
		storage[699] =  11'b10010010000; // [0.5703125]
		storage[700] =  11'b10010001000; // [0.56640625]
		storage[701] =  11'b10010011000; // [0.57421875]
		storage[702] =  11'b10010101000; // [0.58203125]
		storage[703] =  11'b10010110000; // [0.5859375]
		storage[704] =  11'b10010100000; // [0.578125]
		storage[705] =  11'b10001100000; // [0.546875]
		storage[706] =  11'b01110000000; // [0.4375]
		storage[707] =  11'b01001000000; // [0.28125]
		storage[708] =  11'b00110111000; // [0.21484375]
		storage[709] =  11'b00110101000; // [0.20703125]
		storage[710] =  11'b00110110000; // [0.2109375]
		storage[711] =  11'b00111100000; // [0.234375]
		storage[712] =  11'b01001000000; // [0.28125]
		storage[713] =  11'b01100100000; // [0.390625]
		storage[714] =  11'b10000100000; // [0.515625]
		storage[715] =  11'b10011000000; // [0.59375]
		storage[716] =  11'b10011100000; // [0.609375]
		storage[717] =  11'b10011100000; // [0.609375]
		storage[718] =  11'b10011100000; // [0.609375]
		storage[719] =  11'b10011011000; // [0.60546875]
		storage[720] =  11'b10011011000; // [0.60546875]
		storage[721] =  11'b10011010000; // [0.6015625]
		storage[722] =  11'b10011001000; // [0.59765625]
		storage[723] =  11'b10010111000; // [0.58984375]
		storage[724] =  11'b10010101000; // [0.58203125]
		storage[725] =  11'b10010100000; // [0.578125]
		storage[726] =  11'b10010011000; // [0.57421875]
		storage[727] =  11'b10010000000; // [0.5625]
		storage[728] =  11'b10001111000; // [0.55859375]
		storage[729] =  11'b10010010000; // [0.5703125]
		storage[730] =  11'b10010011000; // [0.57421875]
		storage[731] =  11'b10010100000; // [0.578125]
		storage[732] =  11'b10010101000; // [0.58203125]
		storage[733] =  11'b10010100000; // [0.578125]
		storage[734] =  11'b10001100000; // [0.546875]
		storage[735] =  11'b01110111000; // [0.46484375]
		storage[736] =  11'b01011010000; // [0.3515625]
		storage[737] =  11'b01001010000; // [0.2890625]
		storage[738] =  11'b01001111000; // [0.30859375]
		storage[739] =  11'b01100101000; // [0.39453125]
		storage[740] =  11'b10000001000; // [0.50390625]
		storage[741] =  11'b10010011000; // [0.57421875]
		storage[742] =  11'b10011011000; // [0.60546875]
		storage[743] =  11'b10011100000; // [0.609375]
		storage[744] =  11'b10011011000; // [0.60546875]
		storage[745] =  11'b10011011000; // [0.60546875]
		storage[746] =  11'b10011010000; // [0.6015625]
		storage[747] =  11'b10011010000; // [0.6015625]
		storage[748] =  11'b10011010000; // [0.6015625]
		storage[749] =  11'b10011001000; // [0.59765625]
		storage[750] =  11'b10010111000; // [0.58984375]
		storage[751] =  11'b10010101000; // [0.58203125]
		storage[752] =  11'b10010100000; // [0.578125]
		storage[753] =  11'b10010011000; // [0.57421875]
		storage[754] =  11'b10010001000; // [0.56640625]
		storage[755] =  11'b10001110000; // [0.5546875]
		storage[756] =  11'b10001101000; // [0.55078125]
		storage[757] =  11'b10001111000; // [0.55859375]
		storage[758] =  11'b10010010000; // [0.5703125]
		storage[759] =  11'b10010100000; // [0.578125]
		storage[760] =  11'b10010110000; // [0.5859375]
		storage[761] =  11'b10010111000; // [0.58984375]
		storage[762] =  11'b10011000000; // [0.59375]
		storage[763] =  11'b10010100000; // [0.578125]
		storage[764] =  11'b10001100000; // [0.546875]
		storage[765] =  11'b10000110000; // [0.5234375]
		storage[766] =  11'b10001010000; // [0.5390625]
		storage[767] =  11'b10010100000; // [0.578125]
		storage[768] =  11'b10011010000; // [0.6015625]
		storage[769] =  11'b10011100000; // [0.609375]
		storage[770] =  11'b10011100000; // [0.609375]
		storage[771] =  11'b10011011000; // [0.60546875]
		storage[772] =  11'b10011010000; // [0.6015625]
		storage[773] =  11'b10011001000; // [0.59765625]
		storage[774] =  11'b10011001000; // [0.59765625]
		storage[775] =  11'b10011001000; // [0.59765625]
		storage[776] =  11'b10011000000; // [0.59375]
		storage[777] =  11'b10010111000; // [0.58984375]
		storage[778] =  11'b10010101000; // [0.58203125]
		storage[779] =  11'b10010100000; // [0.578125]
		storage[780] =  11'b10010011000; // [0.57421875]
		storage[781] =  11'b10010010000; // [0.5703125]
		storage[782] =  11'b10010000000; // [0.5625]
		storage[783] =  11'b10001101000; // [0.55078125]
	end
endmodule